module sup1v8_n1 (
);

endmodule
