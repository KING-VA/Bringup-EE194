module backingscratchpad_ext(
  input  [12:0] RW0_addr,
  input         RW0_clk,
  input  [63:0] RW0_wdata,
  output [63:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input  [7:0]  RW0_wmask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [11:0] mem_0_0_adr;
  wire  mem_0_0_clk;
  wire [63:0] mem_0_0_din;
  wire [63:0] mem_0_0_q;
  wire  mem_0_0_ren;
  wire  mem_0_0_wen;
  wire [63:0] mem_0_0_wbeb;
  wire  mem_0_0_mcen;
  wire [2:0] mem_0_0_mc;
  wire [1:0] mem_0_0_wa;
  wire [1:0] mem_0_0_wpulse;
  wire  mem_0_0_wpulseen;
  wire  mem_0_0_fwen;
  wire  mem_0_0_clkbyp;
  wire [11:0] mem_1_0_adr;
  wire  mem_1_0_clk;
  wire [63:0] mem_1_0_din;
  wire [63:0] mem_1_0_q;
  wire  mem_1_0_ren;
  wire  mem_1_0_wen;
  wire [63:0] mem_1_0_wbeb;
  wire  mem_1_0_mcen;
  wire [2:0] mem_1_0_mc;
  wire [1:0] mem_1_0_wa;
  wire [1:0] mem_1_0_wpulse;
  wire  mem_1_0_wpulseen;
  wire  mem_1_0_fwen;
  wire  mem_1_0_clkbyp;
  wire  RW0_addr_sel = RW0_addr[12];
  reg  RW0_addr_sel_reg;
  wire [63:0] RW0_rdata_0_0 = mem_0_0_q;
  wire [63:0] RW0_rdata_0 = RW0_rdata_0_0;
  wire [63:0] RW0_rdata_1_0 = mem_1_0_q;
  wire [63:0] RW0_rdata_1 = RW0_rdata_1_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode & RW0_en;
  wire  _GEN_2 = ~RW0_addr_sel;
  wire  _GEN_3 = RW0_wmode & RW0_en;
  wire  _GEN_4 = ~RW0_addr_sel;
  wire  _GEN_5 = RW0_wmask[0];
  wire  _GEN_6 = RW0_wmask[0];
  wire  _GEN_7 = RW0_wmask[0];
  wire [1:0] _GEN_8 = {RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_9 = RW0_wmask[0];
  wire [2:0] _GEN_10 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_11 = RW0_wmask[0];
  wire [3:0] _GEN_12 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_13 = RW0_wmask[0];
  wire [4:0] _GEN_14 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_15 = RW0_wmask[0];
  wire [5:0] _GEN_16 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_17 = RW0_wmask[0];
  wire [6:0] _GEN_18 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_19 = RW0_wmask[1];
  wire [7:0] _GEN_20 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0]};
  wire  _GEN_21 = RW0_wmask[1];
  wire [8:0] _GEN_22 = {RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_23 = RW0_wmask[1];
  wire [9:0] _GEN_24 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_25 = RW0_wmask[1];
  wire [10:0] _GEN_26 = {RW0_wmask[1],_GEN_24};
  wire  _GEN_27 = RW0_wmask[1];
  wire [11:0] _GEN_28 = {RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_29 = RW0_wmask[1];
  wire [12:0] _GEN_30 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_31 = RW0_wmask[1];
  wire [13:0] _GEN_32 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_33 = RW0_wmask[1];
  wire [14:0] _GEN_34 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_35 = RW0_wmask[2];
  wire [15:0] _GEN_36 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_37 = RW0_wmask[2];
  wire [16:0] _GEN_38 = {RW0_wmask[2],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    _GEN_24};
  wire  _GEN_39 = RW0_wmask[2];
  wire [17:0] _GEN_40 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],_GEN_24};
  wire  _GEN_41 = RW0_wmask[2];
  wire [18:0] _GEN_42 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_43 = RW0_wmask[2];
  wire [19:0] _GEN_44 = {RW0_wmask[2],_GEN_42};
  wire  _GEN_45 = RW0_wmask[2];
  wire [20:0] _GEN_46 = {RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_47 = RW0_wmask[2];
  wire [21:0] _GEN_48 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_49 = RW0_wmask[2];
  wire [22:0] _GEN_50 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_51 = RW0_wmask[3];
  wire [23:0] _GEN_52 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_53 = RW0_wmask[3];
  wire [24:0] _GEN_54 = {RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_55 = RW0_wmask[3];
  wire [25:0] _GEN_56 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    _GEN_42};
  wire  _GEN_57 = RW0_wmask[3];
  wire [26:0] _GEN_58 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],_GEN_42};
  wire  _GEN_59 = RW0_wmask[3];
  wire [27:0] _GEN_60 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_61 = RW0_wmask[3];
  wire [28:0] _GEN_62 = {RW0_wmask[3],_GEN_60};
  wire  _GEN_63 = RW0_wmask[3];
  wire [29:0] _GEN_64 = {RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_65 = RW0_wmask[3];
  wire [30:0] _GEN_66 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_67 = RW0_wmask[4];
  wire [31:0] _GEN_68 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_69 = RW0_wmask[4];
  wire [32:0] _GEN_70 = {RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_71 = RW0_wmask[4];
  wire [33:0] _GEN_72 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_73 = RW0_wmask[4];
  wire [34:0] _GEN_74 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    _GEN_60};
  wire  _GEN_75 = RW0_wmask[4];
  wire [35:0] _GEN_76 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],_GEN_60};
  wire  _GEN_77 = RW0_wmask[4];
  wire [36:0] _GEN_78 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_79 = RW0_wmask[4];
  wire [37:0] _GEN_80 = {RW0_wmask[4],_GEN_78};
  wire  _GEN_81 = RW0_wmask[4];
  wire [38:0] _GEN_82 = {RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_83 = RW0_wmask[5];
  wire [39:0] _GEN_84 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_85 = RW0_wmask[5];
  wire [40:0] _GEN_86 = {RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_87 = RW0_wmask[5];
  wire [41:0] _GEN_88 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_89 = RW0_wmask[5];
  wire [42:0] _GEN_90 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_91 = RW0_wmask[5];
  wire [43:0] _GEN_92 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],
    _GEN_78};
  wire  _GEN_93 = RW0_wmask[5];
  wire [44:0] _GEN_94 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],
    RW0_wmask[4],_GEN_78};
  wire  _GEN_95 = RW0_wmask[5];
  wire [45:0] _GEN_96 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],
    RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_97 = RW0_wmask[5];
  wire [46:0] _GEN_98 = {RW0_wmask[5],_GEN_96};
  wire  _GEN_99 = RW0_wmask[6];
  wire [47:0] _GEN_100 = {RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_101 = RW0_wmask[6];
  wire [48:0] _GEN_102 = {RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_103 = RW0_wmask[6];
  wire [49:0] _GEN_104 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_105 = RW0_wmask[6];
  wire [50:0] _GEN_106 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_107 = RW0_wmask[6];
  wire [51:0] _GEN_108 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_109 = RW0_wmask[6];
  wire [52:0] _GEN_110 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],
    _GEN_96};
  wire  _GEN_111 = RW0_wmask[6];
  wire [53:0] _GEN_112 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],
    RW0_wmask[5],_GEN_96};
  wire  _GEN_113 = RW0_wmask[6];
  wire [54:0] _GEN_114 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],
    RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_115 = RW0_wmask[7];
  wire [55:0] _GEN_116 = {RW0_wmask[6],_GEN_114};
  wire  _GEN_117 = RW0_wmask[7];
  wire [56:0] _GEN_118 = {RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_119 = RW0_wmask[7];
  wire [57:0] _GEN_120 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_121 = RW0_wmask[7];
  wire [58:0] _GEN_122 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_123 = RW0_wmask[7];
  wire [59:0] _GEN_124 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_125 = RW0_wmask[7];
  wire [60:0] _GEN_126 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_127 = RW0_wmask[7];
  wire [61:0] _GEN_128 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],
    _GEN_114};
  wire  _GEN_129 = RW0_wmask[7];
  wire [62:0] _GEN_130 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],
    RW0_wmask[6],_GEN_114};
  wire [63:0] _GEN_131 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],
    RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_132 = ~RW0_wmode;
  wire  _GEN_133 = ~RW0_wmode & RW0_en;
  wire  _GEN_134 = RW0_wmode & RW0_en;
  wire  _GEN_135 = RW0_wmask[0];
  wire  _GEN_136 = RW0_wmask[0];
  wire  _GEN_137 = RW0_wmask[0];
  wire [1:0] _GEN_138 = {RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_139 = RW0_wmask[0];
  wire [2:0] _GEN_140 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_141 = RW0_wmask[0];
  wire [3:0] _GEN_142 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_143 = RW0_wmask[0];
  wire [4:0] _GEN_144 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_145 = RW0_wmask[0];
  wire [5:0] _GEN_146 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_147 = RW0_wmask[0];
  wire [6:0] _GEN_148 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_149 = RW0_wmask[1];
  wire [7:0] _GEN_150 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0]};
  wire  _GEN_151 = RW0_wmask[1];
  wire [8:0] _GEN_152 = {RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_153 = RW0_wmask[1];
  wire [9:0] _GEN_154 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_155 = RW0_wmask[1];
  wire [10:0] _GEN_156 = {RW0_wmask[1],_GEN_24};
  wire  _GEN_157 = RW0_wmask[1];
  wire [11:0] _GEN_158 = {RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_159 = RW0_wmask[1];
  wire [12:0] _GEN_160 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_161 = RW0_wmask[1];
  wire [13:0] _GEN_162 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_163 = RW0_wmask[1];
  wire [14:0] _GEN_164 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_165 = RW0_wmask[2];
  wire [15:0] _GEN_166 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_167 = RW0_wmask[2];
  wire [16:0] _GEN_168 = {RW0_wmask[2],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    _GEN_24};
  wire  _GEN_169 = RW0_wmask[2];
  wire [17:0] _GEN_170 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],_GEN_24};
  wire  _GEN_171 = RW0_wmask[2];
  wire [18:0] _GEN_172 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_173 = RW0_wmask[2];
  wire [19:0] _GEN_174 = {RW0_wmask[2],_GEN_42};
  wire  _GEN_175 = RW0_wmask[2];
  wire [20:0] _GEN_176 = {RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_177 = RW0_wmask[2];
  wire [21:0] _GEN_178 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_179 = RW0_wmask[2];
  wire [22:0] _GEN_180 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_181 = RW0_wmask[3];
  wire [23:0] _GEN_182 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_183 = RW0_wmask[3];
  wire [24:0] _GEN_184 = {RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_185 = RW0_wmask[3];
  wire [25:0] _GEN_186 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    _GEN_42};
  wire  _GEN_187 = RW0_wmask[3];
  wire [26:0] _GEN_188 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],_GEN_42};
  wire  _GEN_189 = RW0_wmask[3];
  wire [27:0] _GEN_190 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_191 = RW0_wmask[3];
  wire [28:0] _GEN_192 = {RW0_wmask[3],_GEN_60};
  wire  _GEN_193 = RW0_wmask[3];
  wire [29:0] _GEN_194 = {RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_195 = RW0_wmask[3];
  wire [30:0] _GEN_196 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_197 = RW0_wmask[4];
  wire [31:0] _GEN_198 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_199 = RW0_wmask[4];
  wire [32:0] _GEN_200 = {RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_201 = RW0_wmask[4];
  wire [33:0] _GEN_202 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_203 = RW0_wmask[4];
  wire [34:0] _GEN_204 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    _GEN_60};
  wire  _GEN_205 = RW0_wmask[4];
  wire [35:0] _GEN_206 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],_GEN_60};
  wire  _GEN_207 = RW0_wmask[4];
  wire [36:0] _GEN_208 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_209 = RW0_wmask[4];
  wire [37:0] _GEN_210 = {RW0_wmask[4],_GEN_78};
  wire  _GEN_211 = RW0_wmask[4];
  wire [38:0] _GEN_212 = {RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_213 = RW0_wmask[5];
  wire [39:0] _GEN_214 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_215 = RW0_wmask[5];
  wire [40:0] _GEN_216 = {RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_217 = RW0_wmask[5];
  wire [41:0] _GEN_218 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_219 = RW0_wmask[5];
  wire [42:0] _GEN_220 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_221 = RW0_wmask[5];
  wire [43:0] _GEN_222 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],
    _GEN_78};
  wire  _GEN_223 = RW0_wmask[5];
  wire [44:0] _GEN_224 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],
    RW0_wmask[4],_GEN_78};
  wire  _GEN_225 = RW0_wmask[5];
  wire [45:0] _GEN_226 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],
    RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_227 = RW0_wmask[5];
  wire [46:0] _GEN_228 = {RW0_wmask[5],_GEN_96};
  wire  _GEN_229 = RW0_wmask[6];
  wire [47:0] _GEN_230 = {RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_231 = RW0_wmask[6];
  wire [48:0] _GEN_232 = {RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_233 = RW0_wmask[6];
  wire [49:0] _GEN_234 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_235 = RW0_wmask[6];
  wire [50:0] _GEN_236 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_237 = RW0_wmask[6];
  wire [51:0] _GEN_238 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_239 = RW0_wmask[6];
  wire [52:0] _GEN_240 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],
    _GEN_96};
  wire  _GEN_241 = RW0_wmask[6];
  wire [53:0] _GEN_242 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],
    RW0_wmask[5],_GEN_96};
  wire  _GEN_243 = RW0_wmask[6];
  wire [54:0] _GEN_244 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],
    RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_245 = RW0_wmask[7];
  wire [55:0] _GEN_246 = {RW0_wmask[6],_GEN_114};
  wire  _GEN_247 = RW0_wmask[7];
  wire [56:0] _GEN_248 = {RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_249 = RW0_wmask[7];
  wire [57:0] _GEN_250 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_251 = RW0_wmask[7];
  wire [58:0] _GEN_252 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_253 = RW0_wmask[7];
  wire [59:0] _GEN_254 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_255 = RW0_wmask[7];
  wire [60:0] _GEN_256 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_257 = RW0_wmask[7];
  wire [61:0] _GEN_258 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],
    _GEN_114};
  wire  _GEN_259 = RW0_wmask[7];
  wire [62:0] _GEN_260 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],
    RW0_wmask[6],_GEN_114};
  wire [63:0] _GEN_261 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],
    RW0_wmask[7],RW0_wmask[6],_GEN_114};
  ip224uhdlp1p11rf_4096x64m4b2c1s1_t0r0p0d0a1m1h mem_0_0 (
    .adr(mem_0_0_adr),
    .clk(mem_0_0_clk),
    .din(mem_0_0_din),
    .q(mem_0_0_q),
    .ren(mem_0_0_ren),
    .wen(mem_0_0_wen),
    .wbeb(mem_0_0_wbeb),
    .mcen(mem_0_0_mcen),
    .mc(mem_0_0_mc),
    .wa(mem_0_0_wa),
    .wpulse(mem_0_0_wpulse),
    .wpulseen(mem_0_0_wpulseen),
    .fwen(mem_0_0_fwen),
    .clkbyp(mem_0_0_clkbyp)
  );
  ip224uhdlp1p11rf_4096x64m4b2c1s1_t0r0p0d0a1m1h mem_1_0 (
    .adr(mem_1_0_adr),
    .clk(mem_1_0_clk),
    .din(mem_1_0_din),
    .q(mem_1_0_q),
    .ren(mem_1_0_ren),
    .wen(mem_1_0_wen),
    .wbeb(mem_1_0_wbeb),
    .mcen(mem_1_0_mcen),
    .mc(mem_1_0_mc),
    .wa(mem_1_0_wa),
    .wpulse(mem_1_0_wpulse),
    .wpulseen(mem_1_0_wpulseen),
    .fwen(mem_1_0_fwen),
    .clkbyp(mem_1_0_clkbyp)
  );
  assign RW0_rdata = ~RW0_addr_sel_reg ? RW0_rdata_0_0 : RW0_addr_sel_reg ? RW0_rdata_1_0 : 64'h0;
  assign mem_0_0_adr = RW0_addr[11:0];
  assign mem_0_0_clk = RW0_clk;
  assign mem_0_0_din = RW0_wdata;
  assign mem_0_0_ren = ~RW0_wmode & RW0_en & ~RW0_addr_sel;
  assign mem_0_0_wen = RW0_wmode & RW0_en & ~RW0_addr_sel;
  assign mem_0_0_wbeb = ~_GEN_131;
  assign mem_0_0_mcen = 1'h0;
  assign mem_0_0_mc = 3'h0;
  assign mem_0_0_wa = 2'h0;
  assign mem_0_0_wpulse = 2'h0;
  assign mem_0_0_wpulseen = 1'h1;
  assign mem_0_0_fwen = 1'h0;
  assign mem_0_0_clkbyp = 1'h0;
  assign mem_1_0_adr = RW0_addr[11:0];
  assign mem_1_0_clk = RW0_clk;
  assign mem_1_0_din = RW0_wdata;
  assign mem_1_0_ren = ~RW0_wmode & RW0_en & RW0_addr_sel;
  assign mem_1_0_wen = RW0_wmode & RW0_en & RW0_addr_sel;
  assign mem_1_0_wbeb = ~_GEN_131;
  assign mem_1_0_mcen = 1'h0;
  assign mem_1_0_mc = 3'h0;
  assign mem_1_0_wa = 2'h0;
  assign mem_1_0_wpulse = 2'h0;
  assign mem_1_0_wpulseen = 1'h1;
  assign mem_1_0_fwen = 1'h0;
  assign mem_1_0_clkbyp = 1'h0;
  always @(posedge RW0_clk) begin
    if (RW0_en) begin
      RW0_addr_sel_reg <= RW0_addr_sel;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  RW0_addr_sel_reg = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cc_dir_ext(
  input  [6:0]   RW0_addr,
  input          RW0_clk,
  input  [207:0] RW0_wdata,
  output [207:0] RW0_rdata,
  input          RW0_en,
  input          RW0_wmode,
  input  [7:0]   RW0_wmask
);
  wire [8:0] mem_0_0_adr;
  wire  mem_0_0_clk;
  wire [41:0] mem_0_0_din;
  wire [41:0] mem_0_0_q;
  wire  mem_0_0_ren;
  wire  mem_0_0_wen;
  wire [41:0] mem_0_0_wbeb;
  wire  mem_0_0_mcen;
  wire [2:0] mem_0_0_mc;
  wire [1:0] mem_0_0_wa;
  wire [1:0] mem_0_0_wpulse;
  wire  mem_0_0_wpulseen;
  wire  mem_0_0_fwen;
  wire  mem_0_0_clkbyp;
  wire [8:0] mem_0_1_adr;
  wire  mem_0_1_clk;
  wire [41:0] mem_0_1_din;
  wire [41:0] mem_0_1_q;
  wire  mem_0_1_ren;
  wire  mem_0_1_wen;
  wire [41:0] mem_0_1_wbeb;
  wire  mem_0_1_mcen;
  wire [2:0] mem_0_1_mc;
  wire [1:0] mem_0_1_wa;
  wire [1:0] mem_0_1_wpulse;
  wire  mem_0_1_wpulseen;
  wire  mem_0_1_fwen;
  wire  mem_0_1_clkbyp;
  wire [8:0] mem_0_2_adr;
  wire  mem_0_2_clk;
  wire [41:0] mem_0_2_din;
  wire [41:0] mem_0_2_q;
  wire  mem_0_2_ren;
  wire  mem_0_2_wen;
  wire [41:0] mem_0_2_wbeb;
  wire  mem_0_2_mcen;
  wire [2:0] mem_0_2_mc;
  wire [1:0] mem_0_2_wa;
  wire [1:0] mem_0_2_wpulse;
  wire  mem_0_2_wpulseen;
  wire  mem_0_2_fwen;
  wire  mem_0_2_clkbyp;
  wire [8:0] mem_0_3_adr;
  wire  mem_0_3_clk;
  wire [41:0] mem_0_3_din;
  wire [41:0] mem_0_3_q;
  wire  mem_0_3_ren;
  wire  mem_0_3_wen;
  wire [41:0] mem_0_3_wbeb;
  wire  mem_0_3_mcen;
  wire [2:0] mem_0_3_mc;
  wire [1:0] mem_0_3_wa;
  wire [1:0] mem_0_3_wpulse;
  wire  mem_0_3_wpulseen;
  wire  mem_0_3_fwen;
  wire  mem_0_3_clkbyp;
  wire [8:0] mem_0_4_adr;
  wire  mem_0_4_clk;
  wire [41:0] mem_0_4_din;
  wire [41:0] mem_0_4_q;
  wire  mem_0_4_ren;
  wire  mem_0_4_wen;
  wire [41:0] mem_0_4_wbeb;
  wire  mem_0_4_mcen;
  wire [2:0] mem_0_4_mc;
  wire [1:0] mem_0_4_wa;
  wire [1:0] mem_0_4_wpulse;
  wire  mem_0_4_wpulseen;
  wire  mem_0_4_fwen;
  wire  mem_0_4_clkbyp;
  wire [41:0] RW0_rdata_0_0 = mem_0_0_q;
  wire [41:0] RW0_rdata_0_1 = mem_0_1_q;
  wire [41:0] RW0_rdata_0_2 = mem_0_2_q;
  wire [41:0] RW0_rdata_0_3 = mem_0_3_q;
  wire [39:0] RW0_rdata_0_4 = mem_0_4_q[39:0];
  wire [83:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [125:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [167:0] _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [207:0] RW0_rdata_0 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [83:0] _GEN_3 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [125:0] _GEN_4 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [167:0] _GEN_5 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire  _GEN_6 = ~RW0_wmode;
  wire  _GEN_7 = RW0_wmask[0];
  wire  _GEN_8 = RW0_wmask[0];
  wire  _GEN_9 = RW0_wmask[0];
  wire [1:0] _GEN_10 = {RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_11 = RW0_wmask[0];
  wire [2:0] _GEN_12 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_13 = RW0_wmask[0];
  wire [3:0] _GEN_14 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_15 = RW0_wmask[0];
  wire [4:0] _GEN_16 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_17 = RW0_wmask[0];
  wire [5:0] _GEN_18 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_19 = RW0_wmask[0];
  wire [6:0] _GEN_20 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_21 = RW0_wmask[0];
  wire [7:0] _GEN_22 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0]};
  wire  _GEN_23 = RW0_wmask[0];
  wire [8:0] _GEN_24 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_25 = RW0_wmask[0];
  wire [9:0] _GEN_26 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_27 = RW0_wmask[0];
  wire [10:0] _GEN_28 = {RW0_wmask[0],_GEN_26};
  wire  _GEN_29 = RW0_wmask[0];
  wire [11:0] _GEN_30 = {RW0_wmask[0],RW0_wmask[0],_GEN_26};
  wire  _GEN_31 = RW0_wmask[0];
  wire [12:0] _GEN_32 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_26};
  wire  _GEN_33 = RW0_wmask[0];
  wire [13:0] _GEN_34 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_26};
  wire  _GEN_35 = RW0_wmask[0];
  wire [14:0] _GEN_36 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_26};
  wire  _GEN_37 = RW0_wmask[0];
  wire [15:0] _GEN_38 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_26};
  wire  _GEN_39 = RW0_wmask[0];
  wire [16:0] _GEN_40 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    _GEN_26};
  wire  _GEN_41 = RW0_wmask[0];
  wire [17:0] _GEN_42 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],_GEN_26};
  wire  _GEN_43 = RW0_wmask[0];
  wire [18:0] _GEN_44 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0],_GEN_26};
  wire  _GEN_45 = RW0_wmask[0];
  wire [19:0] _GEN_46 = {RW0_wmask[0],_GEN_44};
  wire  _GEN_47 = RW0_wmask[0];
  wire [20:0] _GEN_48 = {RW0_wmask[0],RW0_wmask[0],_GEN_44};
  wire  _GEN_49 = RW0_wmask[0];
  wire [21:0] _GEN_50 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_44};
  wire  _GEN_51 = RW0_wmask[0];
  wire [22:0] _GEN_52 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_44};
  wire  _GEN_53 = RW0_wmask[0];
  wire [23:0] _GEN_54 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_44};
  wire  _GEN_55 = RW0_wmask[0];
  wire [24:0] _GEN_56 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_44};
  wire  _GEN_57 = RW0_wmask[1];
  wire [25:0] _GEN_58 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    _GEN_44};
  wire  _GEN_59 = RW0_wmask[1];
  wire [26:0] _GEN_60 = {RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],_GEN_44};
  wire  _GEN_61 = RW0_wmask[1];
  wire [27:0] _GEN_62 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0],_GEN_44};
  wire  _GEN_63 = RW0_wmask[1];
  wire [28:0] _GEN_64 = {RW0_wmask[1],_GEN_62};
  wire  _GEN_65 = RW0_wmask[1];
  wire [29:0] _GEN_66 = {RW0_wmask[1],RW0_wmask[1],_GEN_62};
  wire  _GEN_67 = RW0_wmask[1];
  wire [30:0] _GEN_68 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_62};
  wire  _GEN_69 = RW0_wmask[1];
  wire [31:0] _GEN_70 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_62};
  wire  _GEN_71 = RW0_wmask[1];
  wire [32:0] _GEN_72 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_62};
  wire  _GEN_73 = RW0_wmask[1];
  wire [33:0] _GEN_74 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_62};
  wire  _GEN_75 = RW0_wmask[1];
  wire [34:0] _GEN_76 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    _GEN_62};
  wire  _GEN_77 = RW0_wmask[1];
  wire [35:0] _GEN_78 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],_GEN_62};
  wire  _GEN_79 = RW0_wmask[1];
  wire [36:0] _GEN_80 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],RW0_wmask[1],_GEN_62};
  wire  _GEN_81 = RW0_wmask[1];
  wire [37:0] _GEN_82 = {RW0_wmask[1],_GEN_80};
  wire  _GEN_83 = RW0_wmask[1];
  wire [38:0] _GEN_84 = {RW0_wmask[1],RW0_wmask[1],_GEN_80};
  wire  _GEN_85 = RW0_wmask[1];
  wire [39:0] _GEN_86 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_80};
  wire  _GEN_87 = RW0_wmask[1];
  wire [40:0] _GEN_88 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_80};
  wire [41:0] _GEN_89 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_80};
  wire  _GEN_90 = ~RW0_wmode;
  wire  _GEN_91 = RW0_wmask[1];
  wire  _GEN_92 = RW0_wmask[1];
  wire  _GEN_93 = RW0_wmask[1];
  wire [1:0] _GEN_94 = {RW0_wmask[1],RW0_wmask[1]};
  wire  _GEN_95 = RW0_wmask[1];
  wire [2:0] _GEN_96 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1]};
  wire  _GEN_97 = RW0_wmask[1];
  wire [3:0] _GEN_98 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1]};
  wire  _GEN_99 = RW0_wmask[1];
  wire [4:0] _GEN_100 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1]};
  wire  _GEN_101 = RW0_wmask[1];
  wire [5:0] _GEN_102 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1]};
  wire  _GEN_103 = RW0_wmask[1];
  wire [6:0] _GEN_104 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1]};
  wire  _GEN_105 = RW0_wmask[1];
  wire [7:0] _GEN_106 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1]};
  wire  _GEN_107 = RW0_wmask[1];
  wire [8:0] _GEN_108 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],RW0_wmask[1]};
  wire  _GEN_109 = RW0_wmask[2];
  wire [9:0] _GEN_110 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],RW0_wmask[1],RW0_wmask[1]};
  wire  _GEN_111 = RW0_wmask[2];
  wire [10:0] _GEN_112 = {RW0_wmask[2],_GEN_110};
  wire  _GEN_113 = RW0_wmask[2];
  wire [11:0] _GEN_114 = {RW0_wmask[2],RW0_wmask[2],_GEN_110};
  wire  _GEN_115 = RW0_wmask[2];
  wire [12:0] _GEN_116 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_110};
  wire  _GEN_117 = RW0_wmask[2];
  wire [13:0] _GEN_118 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_110};
  wire  _GEN_119 = RW0_wmask[2];
  wire [14:0] _GEN_120 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_110};
  wire  _GEN_121 = RW0_wmask[2];
  wire [15:0] _GEN_122 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_110};
  wire  _GEN_123 = RW0_wmask[2];
  wire [16:0] _GEN_124 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    _GEN_110};
  wire  _GEN_125 = RW0_wmask[2];
  wire [17:0] _GEN_126 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],_GEN_110};
  wire  _GEN_127 = RW0_wmask[2];
  wire [18:0] _GEN_128 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],RW0_wmask[2],_GEN_110};
  wire  _GEN_129 = RW0_wmask[2];
  wire [19:0] _GEN_130 = {RW0_wmask[2],_GEN_128};
  wire  _GEN_131 = RW0_wmask[2];
  wire [20:0] _GEN_132 = {RW0_wmask[2],RW0_wmask[2],_GEN_128};
  wire  _GEN_133 = RW0_wmask[2];
  wire [21:0] _GEN_134 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_128};
  wire  _GEN_135 = RW0_wmask[2];
  wire [22:0] _GEN_136 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_128};
  wire  _GEN_137 = RW0_wmask[2];
  wire [23:0] _GEN_138 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_128};
  wire  _GEN_139 = RW0_wmask[2];
  wire [24:0] _GEN_140 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_128};
  wire  _GEN_141 = RW0_wmask[2];
  wire [25:0] _GEN_142 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    _GEN_128};
  wire  _GEN_143 = RW0_wmask[2];
  wire [26:0] _GEN_144 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],_GEN_128};
  wire  _GEN_145 = RW0_wmask[2];
  wire [27:0] _GEN_146 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],RW0_wmask[2],_GEN_128};
  wire  _GEN_147 = RW0_wmask[2];
  wire [28:0] _GEN_148 = {RW0_wmask[2],_GEN_146};
  wire  _GEN_149 = RW0_wmask[2];
  wire [29:0] _GEN_150 = {RW0_wmask[2],RW0_wmask[2],_GEN_146};
  wire  _GEN_151 = RW0_wmask[2];
  wire [30:0] _GEN_152 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_146};
  wire  _GEN_153 = RW0_wmask[2];
  wire [31:0] _GEN_154 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_146};
  wire  _GEN_155 = RW0_wmask[2];
  wire [32:0] _GEN_156 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_146};
  wire  _GEN_157 = RW0_wmask[2];
  wire [33:0] _GEN_158 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_146};
  wire  _GEN_159 = RW0_wmask[2];
  wire [34:0] _GEN_160 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    _GEN_146};
  wire  _GEN_161 = RW0_wmask[3];
  wire [35:0] _GEN_162 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],_GEN_146};
  wire  _GEN_163 = RW0_wmask[3];
  wire [36:0] _GEN_164 = {RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],RW0_wmask[2],_GEN_146};
  wire  _GEN_165 = RW0_wmask[3];
  wire [37:0] _GEN_166 = {RW0_wmask[3],_GEN_164};
  wire  _GEN_167 = RW0_wmask[3];
  wire [38:0] _GEN_168 = {RW0_wmask[3],RW0_wmask[3],_GEN_164};
  wire  _GEN_169 = RW0_wmask[3];
  wire [39:0] _GEN_170 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_164};
  wire  _GEN_171 = RW0_wmask[3];
  wire [40:0] _GEN_172 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_164};
  wire [41:0] _GEN_173 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_164};
  wire  _GEN_174 = ~RW0_wmode;
  wire  _GEN_175 = RW0_wmask[3];
  wire  _GEN_176 = RW0_wmask[3];
  wire  _GEN_177 = RW0_wmask[3];
  wire [1:0] _GEN_178 = {RW0_wmask[3],RW0_wmask[3]};
  wire  _GEN_179 = RW0_wmask[3];
  wire [2:0] _GEN_180 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3]};
  wire  _GEN_181 = RW0_wmask[3];
  wire [3:0] _GEN_182 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3]};
  wire  _GEN_183 = RW0_wmask[3];
  wire [4:0] _GEN_184 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3]};
  wire  _GEN_185 = RW0_wmask[3];
  wire [5:0] _GEN_186 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3]};
  wire  _GEN_187 = RW0_wmask[3];
  wire [6:0] _GEN_188 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3]};
  wire  _GEN_189 = RW0_wmask[3];
  wire [7:0] _GEN_190 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3]};
  wire  _GEN_191 = RW0_wmask[3];
  wire [8:0] _GEN_192 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],RW0_wmask[3]};
  wire  _GEN_193 = RW0_wmask[3];
  wire [9:0] _GEN_194 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],RW0_wmask[3],RW0_wmask[3]};
  wire  _GEN_195 = RW0_wmask[3];
  wire [10:0] _GEN_196 = {RW0_wmask[3],_GEN_194};
  wire  _GEN_197 = RW0_wmask[3];
  wire [11:0] _GEN_198 = {RW0_wmask[3],RW0_wmask[3],_GEN_194};
  wire  _GEN_199 = RW0_wmask[3];
  wire [12:0] _GEN_200 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_194};
  wire  _GEN_201 = RW0_wmask[3];
  wire [13:0] _GEN_202 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_194};
  wire  _GEN_203 = RW0_wmask[3];
  wire [14:0] _GEN_204 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_194};
  wire  _GEN_205 = RW0_wmask[3];
  wire [15:0] _GEN_206 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_194};
  wire  _GEN_207 = RW0_wmask[3];
  wire [16:0] _GEN_208 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    _GEN_194};
  wire  _GEN_209 = RW0_wmask[3];
  wire [17:0] _GEN_210 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],_GEN_194};
  wire  _GEN_211 = RW0_wmask[3];
  wire [18:0] _GEN_212 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],RW0_wmask[3],_GEN_194};
  wire  _GEN_213 = RW0_wmask[4];
  wire [19:0] _GEN_214 = {RW0_wmask[3],_GEN_212};
  wire  _GEN_215 = RW0_wmask[4];
  wire [20:0] _GEN_216 = {RW0_wmask[4],RW0_wmask[3],_GEN_212};
  wire  _GEN_217 = RW0_wmask[4];
  wire [21:0] _GEN_218 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],_GEN_212};
  wire  _GEN_219 = RW0_wmask[4];
  wire [22:0] _GEN_220 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],_GEN_212};
  wire  _GEN_221 = RW0_wmask[4];
  wire [23:0] _GEN_222 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],_GEN_212};
  wire  _GEN_223 = RW0_wmask[4];
  wire [24:0] _GEN_224 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],_GEN_212};
  wire  _GEN_225 = RW0_wmask[4];
  wire [25:0] _GEN_226 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],
    _GEN_212};
  wire  _GEN_227 = RW0_wmask[4];
  wire [26:0] _GEN_228 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],
    RW0_wmask[3],_GEN_212};
  wire  _GEN_229 = RW0_wmask[4];
  wire [27:0] _GEN_230 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],
    RW0_wmask[4],RW0_wmask[3],_GEN_212};
  wire  _GEN_231 = RW0_wmask[4];
  wire [28:0] _GEN_232 = {RW0_wmask[4],_GEN_230};
  wire  _GEN_233 = RW0_wmask[4];
  wire [29:0] _GEN_234 = {RW0_wmask[4],RW0_wmask[4],_GEN_230};
  wire  _GEN_235 = RW0_wmask[4];
  wire [30:0] _GEN_236 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_230};
  wire  _GEN_237 = RW0_wmask[4];
  wire [31:0] _GEN_238 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_230};
  wire  _GEN_239 = RW0_wmask[4];
  wire [32:0] _GEN_240 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_230};
  wire  _GEN_241 = RW0_wmask[4];
  wire [33:0] _GEN_242 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_230};
  wire  _GEN_243 = RW0_wmask[4];
  wire [34:0] _GEN_244 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],
    _GEN_230};
  wire  _GEN_245 = RW0_wmask[4];
  wire [35:0] _GEN_246 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],
    RW0_wmask[4],_GEN_230};
  wire  _GEN_247 = RW0_wmask[4];
  wire [36:0] _GEN_248 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],
    RW0_wmask[4],RW0_wmask[4],_GEN_230};
  wire  _GEN_249 = RW0_wmask[4];
  wire [37:0] _GEN_250 = {RW0_wmask[4],_GEN_248};
  wire  _GEN_251 = RW0_wmask[4];
  wire [38:0] _GEN_252 = {RW0_wmask[4],RW0_wmask[4],_GEN_248};
  wire  _GEN_253 = RW0_wmask[4];
  wire [39:0] _GEN_254 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_248};
  wire  _GEN_255 = RW0_wmask[4];
  wire [40:0] _GEN_256 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_248};
  wire [41:0] _GEN_257 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_248};
  wire  _GEN_258 = ~RW0_wmode;
  wire  _GEN_259 = RW0_wmask[4];
  wire  _GEN_260 = RW0_wmask[4];
  wire  _GEN_261 = RW0_wmask[4];
  wire [1:0] _GEN_262 = {RW0_wmask[4],RW0_wmask[4]};
  wire  _GEN_263 = RW0_wmask[4];
  wire [2:0] _GEN_264 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4]};
  wire  _GEN_265 = RW0_wmask[5];
  wire [3:0] _GEN_266 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4]};
  wire  _GEN_267 = RW0_wmask[5];
  wire [4:0] _GEN_268 = {RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4]};
  wire  _GEN_269 = RW0_wmask[5];
  wire [5:0] _GEN_270 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4]};
  wire  _GEN_271 = RW0_wmask[5];
  wire [6:0] _GEN_272 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4]};
  wire  _GEN_273 = RW0_wmask[5];
  wire [7:0] _GEN_274 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],
    RW0_wmask[4]};
  wire  _GEN_275 = RW0_wmask[5];
  wire [8:0] _GEN_276 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],
    RW0_wmask[4],RW0_wmask[4]};
  wire  _GEN_277 = RW0_wmask[5];
  wire [9:0] _GEN_278 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],
    RW0_wmask[4],RW0_wmask[4],RW0_wmask[4]};
  wire  _GEN_279 = RW0_wmask[5];
  wire [10:0] _GEN_280 = {RW0_wmask[5],_GEN_278};
  wire  _GEN_281 = RW0_wmask[5];
  wire [11:0] _GEN_282 = {RW0_wmask[5],RW0_wmask[5],_GEN_278};
  wire  _GEN_283 = RW0_wmask[5];
  wire [12:0] _GEN_284 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],_GEN_278};
  wire  _GEN_285 = RW0_wmask[5];
  wire [13:0] _GEN_286 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],_GEN_278};
  wire  _GEN_287 = RW0_wmask[5];
  wire [14:0] _GEN_288 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],_GEN_278};
  wire  _GEN_289 = RW0_wmask[5];
  wire [15:0] _GEN_290 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],_GEN_278};
  wire  _GEN_291 = RW0_wmask[5];
  wire [16:0] _GEN_292 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],
    _GEN_278};
  wire  _GEN_293 = RW0_wmask[5];
  wire [17:0] _GEN_294 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],
    RW0_wmask[5],_GEN_278};
  wire  _GEN_295 = RW0_wmask[5];
  wire [18:0] _GEN_296 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],
    RW0_wmask[5],RW0_wmask[5],_GEN_278};
  wire  _GEN_297 = RW0_wmask[5];
  wire [19:0] _GEN_298 = {RW0_wmask[5],_GEN_296};
  wire  _GEN_299 = RW0_wmask[5];
  wire [20:0] _GEN_300 = {RW0_wmask[5],RW0_wmask[5],_GEN_296};
  wire  _GEN_301 = RW0_wmask[5];
  wire [21:0] _GEN_302 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],_GEN_296};
  wire  _GEN_303 = RW0_wmask[5];
  wire [22:0] _GEN_304 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],_GEN_296};
  wire  _GEN_305 = RW0_wmask[5];
  wire [23:0] _GEN_306 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],_GEN_296};
  wire  _GEN_307 = RW0_wmask[5];
  wire [24:0] _GEN_308 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],_GEN_296};
  wire  _GEN_309 = RW0_wmask[5];
  wire [25:0] _GEN_310 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],
    _GEN_296};
  wire  _GEN_311 = RW0_wmask[5];
  wire [26:0] _GEN_312 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],
    RW0_wmask[5],_GEN_296};
  wire  _GEN_313 = RW0_wmask[5];
  wire [27:0] _GEN_314 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],
    RW0_wmask[5],RW0_wmask[5],_GEN_296};
  wire  _GEN_315 = RW0_wmask[5];
  wire [28:0] _GEN_316 = {RW0_wmask[5],_GEN_314};
  wire  _GEN_317 = RW0_wmask[6];
  wire [29:0] _GEN_318 = {RW0_wmask[5],RW0_wmask[5],_GEN_314};
  wire  _GEN_319 = RW0_wmask[6];
  wire [30:0] _GEN_320 = {RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_314};
  wire  _GEN_321 = RW0_wmask[6];
  wire [31:0] _GEN_322 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_314};
  wire  _GEN_323 = RW0_wmask[6];
  wire [32:0] _GEN_324 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_314};
  wire  _GEN_325 = RW0_wmask[6];
  wire [33:0] _GEN_326 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_314};
  wire  _GEN_327 = RW0_wmask[6];
  wire [34:0] _GEN_328 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],
    _GEN_314};
  wire  _GEN_329 = RW0_wmask[6];
  wire [35:0] _GEN_330 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],
    RW0_wmask[5],_GEN_314};
  wire  _GEN_331 = RW0_wmask[6];
  wire [36:0] _GEN_332 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],
    RW0_wmask[5],RW0_wmask[5],_GEN_314};
  wire  _GEN_333 = RW0_wmask[6];
  wire [37:0] _GEN_334 = {RW0_wmask[6],_GEN_332};
  wire  _GEN_335 = RW0_wmask[6];
  wire [38:0] _GEN_336 = {RW0_wmask[6],RW0_wmask[6],_GEN_332};
  wire  _GEN_337 = RW0_wmask[6];
  wire [39:0] _GEN_338 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],_GEN_332};
  wire  _GEN_339 = RW0_wmask[6];
  wire [40:0] _GEN_340 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],_GEN_332};
  wire [41:0] _GEN_341 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],_GEN_332};
  wire [39:0] _GEN_342 = RW0_wdata[207:168];
  wire  _GEN_343 = ~RW0_wmode;
  wire  _GEN_344 = RW0_wmask[6];
  wire  _GEN_345 = RW0_wmask[6];
  wire  _GEN_346 = RW0_wmask[6];
  wire [1:0] _GEN_347 = {RW0_wmask[6],RW0_wmask[6]};
  wire  _GEN_348 = RW0_wmask[6];
  wire [2:0] _GEN_349 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6]};
  wire  _GEN_350 = RW0_wmask[6];
  wire [3:0] _GEN_351 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6]};
  wire  _GEN_352 = RW0_wmask[6];
  wire [4:0] _GEN_353 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6]};
  wire  _GEN_354 = RW0_wmask[6];
  wire [5:0] _GEN_355 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6]};
  wire  _GEN_356 = RW0_wmask[6];
  wire [6:0] _GEN_357 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6]};
  wire  _GEN_358 = RW0_wmask[6];
  wire [7:0] _GEN_359 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],
    RW0_wmask[6]};
  wire  _GEN_360 = RW0_wmask[6];
  wire [8:0] _GEN_361 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],
    RW0_wmask[6],RW0_wmask[6]};
  wire  _GEN_362 = RW0_wmask[6];
  wire [9:0] _GEN_363 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],
    RW0_wmask[6],RW0_wmask[6],RW0_wmask[6]};
  wire  _GEN_364 = RW0_wmask[6];
  wire [10:0] _GEN_365 = {RW0_wmask[6],_GEN_363};
  wire  _GEN_366 = RW0_wmask[6];
  wire [11:0] _GEN_367 = {RW0_wmask[6],RW0_wmask[6],_GEN_363};
  wire  _GEN_368 = RW0_wmask[6];
  wire [12:0] _GEN_369 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],_GEN_363};
  wire  _GEN_370 = RW0_wmask[7];
  wire [13:0] _GEN_371 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],_GEN_363};
  wire  _GEN_372 = RW0_wmask[7];
  wire [14:0] _GEN_373 = {RW0_wmask[7],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],_GEN_363};
  wire  _GEN_374 = RW0_wmask[7];
  wire [15:0] _GEN_375 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],_GEN_363};
  wire  _GEN_376 = RW0_wmask[7];
  wire [16:0] _GEN_377 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],
    _GEN_363};
  wire  _GEN_378 = RW0_wmask[7];
  wire [17:0] _GEN_379 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],
    RW0_wmask[6],_GEN_363};
  wire  _GEN_380 = RW0_wmask[7];
  wire [18:0] _GEN_381 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],RW0_wmask[6],
    RW0_wmask[6],RW0_wmask[6],_GEN_363};
  wire  _GEN_382 = RW0_wmask[7];
  wire [19:0] _GEN_383 = {RW0_wmask[7],_GEN_381};
  wire  _GEN_384 = RW0_wmask[7];
  wire [20:0] _GEN_385 = {RW0_wmask[7],RW0_wmask[7],_GEN_381};
  wire  _GEN_386 = RW0_wmask[7];
  wire [21:0] _GEN_387 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],_GEN_381};
  wire  _GEN_388 = RW0_wmask[7];
  wire [22:0] _GEN_389 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],_GEN_381};
  wire  _GEN_390 = RW0_wmask[7];
  wire [23:0] _GEN_391 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],_GEN_381};
  wire  _GEN_392 = RW0_wmask[7];
  wire [24:0] _GEN_393 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],_GEN_381};
  wire  _GEN_394 = RW0_wmask[7];
  wire [25:0] _GEN_395 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],
    _GEN_381};
  wire  _GEN_396 = RW0_wmask[7];
  wire [26:0] _GEN_397 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],
    RW0_wmask[7],_GEN_381};
  wire  _GEN_398 = RW0_wmask[7];
  wire [27:0] _GEN_399 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],
    RW0_wmask[7],RW0_wmask[7],_GEN_381};
  wire  _GEN_400 = RW0_wmask[7];
  wire [28:0] _GEN_401 = {RW0_wmask[7],_GEN_399};
  wire  _GEN_402 = RW0_wmask[7];
  wire [29:0] _GEN_403 = {RW0_wmask[7],RW0_wmask[7],_GEN_399};
  wire  _GEN_404 = RW0_wmask[7];
  wire [30:0] _GEN_405 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],_GEN_399};
  wire  _GEN_406 = RW0_wmask[7];
  wire [31:0] _GEN_407 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],_GEN_399};
  wire  _GEN_408 = RW0_wmask[7];
  wire [32:0] _GEN_409 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],_GEN_399};
  wire  _GEN_410 = RW0_wmask[7];
  wire [33:0] _GEN_411 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],_GEN_399};
  wire  _GEN_412 = RW0_wmask[7];
  wire [34:0] _GEN_413 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],
    _GEN_399};
  wire  _GEN_414 = RW0_wmask[7];
  wire [35:0] _GEN_415 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],
    RW0_wmask[7],_GEN_399};
  wire  _GEN_416 = RW0_wmask[7];
  wire [36:0] _GEN_417 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],
    RW0_wmask[7],RW0_wmask[7],_GEN_399};
  wire  _GEN_418 = RW0_wmask[7];
  wire [37:0] _GEN_419 = {RW0_wmask[7],_GEN_417};
  wire  _GEN_420 = RW0_wmask[7];
  wire [38:0] _GEN_421 = {RW0_wmask[7],RW0_wmask[7],_GEN_417};
  wire [39:0] _GEN_422 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],_GEN_417};
  wire [40:0] _GEN_423 = {1'h0,RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],_GEN_417};
  wire [41:0] _GEN_424 = {1'h0,1'h0,RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],_GEN_417};
  ip224uhdlp1p11rf_512x42m4b2c1s1_t0r0p0d0a1m1h mem_0_0 (
    .adr(mem_0_0_adr),
    .clk(mem_0_0_clk),
    .din(mem_0_0_din),
    .q(mem_0_0_q),
    .ren(mem_0_0_ren),
    .wen(mem_0_0_wen),
    .wbeb(mem_0_0_wbeb),
    .mcen(mem_0_0_mcen),
    .mc(mem_0_0_mc),
    .wa(mem_0_0_wa),
    .wpulse(mem_0_0_wpulse),
    .wpulseen(mem_0_0_wpulseen),
    .fwen(mem_0_0_fwen),
    .clkbyp(mem_0_0_clkbyp)
  );
  ip224uhdlp1p11rf_512x42m4b2c1s1_t0r0p0d0a1m1h mem_0_1 (
    .adr(mem_0_1_adr),
    .clk(mem_0_1_clk),
    .din(mem_0_1_din),
    .q(mem_0_1_q),
    .ren(mem_0_1_ren),
    .wen(mem_0_1_wen),
    .wbeb(mem_0_1_wbeb),
    .mcen(mem_0_1_mcen),
    .mc(mem_0_1_mc),
    .wa(mem_0_1_wa),
    .wpulse(mem_0_1_wpulse),
    .wpulseen(mem_0_1_wpulseen),
    .fwen(mem_0_1_fwen),
    .clkbyp(mem_0_1_clkbyp)
  );
  ip224uhdlp1p11rf_512x42m4b2c1s1_t0r0p0d0a1m1h mem_0_2 (
    .adr(mem_0_2_adr),
    .clk(mem_0_2_clk),
    .din(mem_0_2_din),
    .q(mem_0_2_q),
    .ren(mem_0_2_ren),
    .wen(mem_0_2_wen),
    .wbeb(mem_0_2_wbeb),
    .mcen(mem_0_2_mcen),
    .mc(mem_0_2_mc),
    .wa(mem_0_2_wa),
    .wpulse(mem_0_2_wpulse),
    .wpulseen(mem_0_2_wpulseen),
    .fwen(mem_0_2_fwen),
    .clkbyp(mem_0_2_clkbyp)
  );
  ip224uhdlp1p11rf_512x42m4b2c1s1_t0r0p0d0a1m1h mem_0_3 (
    .adr(mem_0_3_adr),
    .clk(mem_0_3_clk),
    .din(mem_0_3_din),
    .q(mem_0_3_q),
    .ren(mem_0_3_ren),
    .wen(mem_0_3_wen),
    .wbeb(mem_0_3_wbeb),
    .mcen(mem_0_3_mcen),
    .mc(mem_0_3_mc),
    .wa(mem_0_3_wa),
    .wpulse(mem_0_3_wpulse),
    .wpulseen(mem_0_3_wpulseen),
    .fwen(mem_0_3_fwen),
    .clkbyp(mem_0_3_clkbyp)
  );
  ip224uhdlp1p11rf_512x42m4b2c1s1_t0r0p0d0a1m1h mem_0_4 (
    .adr(mem_0_4_adr),
    .clk(mem_0_4_clk),
    .din(mem_0_4_din),
    .q(mem_0_4_q),
    .ren(mem_0_4_ren),
    .wen(mem_0_4_wen),
    .wbeb(mem_0_4_wbeb),
    .mcen(mem_0_4_mcen),
    .mc(mem_0_4_mc),
    .wa(mem_0_4_wa),
    .wpulse(mem_0_4_wpulse),
    .wpulseen(mem_0_4_wpulseen),
    .fwen(mem_0_4_fwen),
    .clkbyp(mem_0_4_clkbyp)
  );
  assign RW0_rdata = {RW0_rdata_0_4,_GEN_2};
  assign mem_0_0_adr = {{2'd0}, RW0_addr};
  assign mem_0_0_clk = RW0_clk;
  assign mem_0_0_din = RW0_wdata[41:0];
  assign mem_0_0_ren = ~RW0_wmode & RW0_en;
  assign mem_0_0_wen = RW0_wmode & RW0_en;
  assign mem_0_0_wbeb = ~_GEN_89;
  assign mem_0_0_mcen = 1'h0;
  assign mem_0_0_mc = 3'h0;
  assign mem_0_0_wa = 2'h0;
  assign mem_0_0_wpulse = 2'h0;
  assign mem_0_0_wpulseen = 1'h1;
  assign mem_0_0_fwen = 1'h0;
  assign mem_0_0_clkbyp = 1'h0;
  assign mem_0_1_adr = {{2'd0}, RW0_addr};
  assign mem_0_1_clk = RW0_clk;
  assign mem_0_1_din = RW0_wdata[83:42];
  assign mem_0_1_ren = ~RW0_wmode & RW0_en;
  assign mem_0_1_wen = RW0_wmode & RW0_en;
  assign mem_0_1_wbeb = ~_GEN_173;
  assign mem_0_1_mcen = 1'h0;
  assign mem_0_1_mc = 3'h0;
  assign mem_0_1_wa = 2'h0;
  assign mem_0_1_wpulse = 2'h0;
  assign mem_0_1_wpulseen = 1'h1;
  assign mem_0_1_fwen = 1'h0;
  assign mem_0_1_clkbyp = 1'h0;
  assign mem_0_2_adr = {{2'd0}, RW0_addr};
  assign mem_0_2_clk = RW0_clk;
  assign mem_0_2_din = RW0_wdata[125:84];
  assign mem_0_2_ren = ~RW0_wmode & RW0_en;
  assign mem_0_2_wen = RW0_wmode & RW0_en;
  assign mem_0_2_wbeb = ~_GEN_257;
  assign mem_0_2_mcen = 1'h0;
  assign mem_0_2_mc = 3'h0;
  assign mem_0_2_wa = 2'h0;
  assign mem_0_2_wpulse = 2'h0;
  assign mem_0_2_wpulseen = 1'h1;
  assign mem_0_2_fwen = 1'h0;
  assign mem_0_2_clkbyp = 1'h0;
  assign mem_0_3_adr = {{2'd0}, RW0_addr};
  assign mem_0_3_clk = RW0_clk;
  assign mem_0_3_din = RW0_wdata[167:126];
  assign mem_0_3_ren = ~RW0_wmode & RW0_en;
  assign mem_0_3_wen = RW0_wmode & RW0_en;
  assign mem_0_3_wbeb = ~_GEN_341;
  assign mem_0_3_mcen = 1'h0;
  assign mem_0_3_mc = 3'h0;
  assign mem_0_3_wa = 2'h0;
  assign mem_0_3_wpulse = 2'h0;
  assign mem_0_3_wpulseen = 1'h1;
  assign mem_0_3_fwen = 1'h0;
  assign mem_0_3_clkbyp = 1'h0;
  assign mem_0_4_adr = {{2'd0}, RW0_addr};
  assign mem_0_4_clk = RW0_clk;
  assign mem_0_4_din = {{2'd0}, RW0_wdata[207:168]};
  assign mem_0_4_ren = ~RW0_wmode & RW0_en;
  assign mem_0_4_wen = RW0_wmode & RW0_en;
  assign mem_0_4_wbeb = ~_GEN_424;
  assign mem_0_4_mcen = 1'h0;
  assign mem_0_4_mc = 3'h0;
  assign mem_0_4_wa = 2'h0;
  assign mem_0_4_wpulse = 2'h0;
  assign mem_0_4_wpulseen = 1'h1;
  assign mem_0_4_fwen = 1'h0;
  assign mem_0_4_clkbyp = 1'h0;
endmodule
module cc_banks_0_ext(
  input  [10:0] RW0_addr,
  input         RW0_clk,
  input  [63:0] RW0_wdata,
  output [63:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [9:0] mem_0_0_adr;
  wire  mem_0_0_clk;
  wire [63:0] mem_0_0_din;
  wire [63:0] mem_0_0_q;
  wire  mem_0_0_ren;
  wire  mem_0_0_wen;
  wire [63:0] mem_0_0_wbeb;
  wire  mem_0_0_mcen;
  wire [2:0] mem_0_0_mc;
  wire [1:0] mem_0_0_wa;
  wire [1:0] mem_0_0_wpulse;
  wire  mem_0_0_wpulseen;
  wire  mem_0_0_fwen;
  wire  mem_0_0_clkbyp;
  wire [9:0] mem_1_0_adr;
  wire  mem_1_0_clk;
  wire [63:0] mem_1_0_din;
  wire [63:0] mem_1_0_q;
  wire  mem_1_0_ren;
  wire  mem_1_0_wen;
  wire [63:0] mem_1_0_wbeb;
  wire  mem_1_0_mcen;
  wire [2:0] mem_1_0_mc;
  wire [1:0] mem_1_0_wa;
  wire [1:0] mem_1_0_wpulse;
  wire  mem_1_0_wpulseen;
  wire  mem_1_0_fwen;
  wire  mem_1_0_clkbyp;
  wire  RW0_addr_sel = RW0_addr[10];
  reg  RW0_addr_sel_reg;
  wire [63:0] RW0_rdata_0_0 = mem_0_0_q;
  wire [63:0] RW0_rdata_0 = RW0_rdata_0_0;
  wire [63:0] RW0_rdata_1_0 = mem_1_0_q;
  wire [63:0] RW0_rdata_1 = RW0_rdata_1_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode & RW0_en;
  wire  _GEN_2 = ~RW0_addr_sel;
  wire  _GEN_3 = RW0_wmode & RW0_en;
  wire  _GEN_4 = ~RW0_addr_sel;
  wire  _GEN_5 = ~RW0_wmode;
  wire  _GEN_6 = ~RW0_wmode & RW0_en;
  wire  _GEN_7 = RW0_wmode & RW0_en;
  ip224uhdlp1p11rf_1024x64m4b2c1s1_t0r0p0d0a1m1h mem_0_0 (
    .adr(mem_0_0_adr),
    .clk(mem_0_0_clk),
    .din(mem_0_0_din),
    .q(mem_0_0_q),
    .ren(mem_0_0_ren),
    .wen(mem_0_0_wen),
    .wbeb(mem_0_0_wbeb),
    .mcen(mem_0_0_mcen),
    .mc(mem_0_0_mc),
    .wa(mem_0_0_wa),
    .wpulse(mem_0_0_wpulse),
    .wpulseen(mem_0_0_wpulseen),
    .fwen(mem_0_0_fwen),
    .clkbyp(mem_0_0_clkbyp)
  );
  ip224uhdlp1p11rf_1024x64m4b2c1s1_t0r0p0d0a1m1h mem_1_0 (
    .adr(mem_1_0_adr),
    .clk(mem_1_0_clk),
    .din(mem_1_0_din),
    .q(mem_1_0_q),
    .ren(mem_1_0_ren),
    .wen(mem_1_0_wen),
    .wbeb(mem_1_0_wbeb),
    .mcen(mem_1_0_mcen),
    .mc(mem_1_0_mc),
    .wa(mem_1_0_wa),
    .wpulse(mem_1_0_wpulse),
    .wpulseen(mem_1_0_wpulseen),
    .fwen(mem_1_0_fwen),
    .clkbyp(mem_1_0_clkbyp)
  );
  assign RW0_rdata = ~RW0_addr_sel_reg ? RW0_rdata_0_0 : RW0_addr_sel_reg ? RW0_rdata_1_0 : 64'h0;
  assign mem_0_0_adr = RW0_addr[9:0];
  assign mem_0_0_clk = RW0_clk;
  assign mem_0_0_din = RW0_wdata;
  assign mem_0_0_ren = ~RW0_wmode & RW0_en & ~RW0_addr_sel;
  assign mem_0_0_wen = RW0_wmode & RW0_en & ~RW0_addr_sel;
  assign mem_0_0_wbeb = 64'h0;
  assign mem_0_0_mcen = 1'h0;
  assign mem_0_0_mc = 3'h0;
  assign mem_0_0_wa = 2'h0;
  assign mem_0_0_wpulse = 2'h0;
  assign mem_0_0_wpulseen = 1'h1;
  assign mem_0_0_fwen = 1'h0;
  assign mem_0_0_clkbyp = 1'h0;
  assign mem_1_0_adr = RW0_addr[9:0];
  assign mem_1_0_clk = RW0_clk;
  assign mem_1_0_din = RW0_wdata;
  assign mem_1_0_ren = ~RW0_wmode & RW0_en & RW0_addr_sel;
  assign mem_1_0_wen = RW0_wmode & RW0_en & RW0_addr_sel;
  assign mem_1_0_wbeb = 64'h0;
  assign mem_1_0_mcen = 1'h0;
  assign mem_1_0_mc = 3'h0;
  assign mem_1_0_wa = 2'h0;
  assign mem_1_0_wpulse = 2'h0;
  assign mem_1_0_wpulseen = 1'h1;
  assign mem_1_0_fwen = 1'h0;
  assign mem_1_0_clkbyp = 1'h0;
  always @(posedge RW0_clk) begin
    if (RW0_en) begin
      RW0_addr_sel_reg <= RW0_addr_sel;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  RW0_addr_sel_reg = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module data_arrays_0_ext(
  input  [8:0]   RW0_addr,
  input          RW0_clk,
  input  [255:0] RW0_wdata,
  output [255:0] RW0_rdata,
  input          RW0_en,
  input          RW0_wmode,
  input  [31:0]  RW0_wmask
);
  wire [8:0] mem_0_0_adr;
  wire  mem_0_0_clk;
  wire [63:0] mem_0_0_din;
  wire [63:0] mem_0_0_q;
  wire  mem_0_0_ren;
  wire  mem_0_0_wen;
  wire [63:0] mem_0_0_wbeb;
  wire  mem_0_0_mcen;
  wire [2:0] mem_0_0_mc;
  wire [1:0] mem_0_0_wa;
  wire [1:0] mem_0_0_wpulse;
  wire  mem_0_0_wpulseen;
  wire  mem_0_0_fwen;
  wire  mem_0_0_clkbyp;
  wire [8:0] mem_0_1_adr;
  wire  mem_0_1_clk;
  wire [63:0] mem_0_1_din;
  wire [63:0] mem_0_1_q;
  wire  mem_0_1_ren;
  wire  mem_0_1_wen;
  wire [63:0] mem_0_1_wbeb;
  wire  mem_0_1_mcen;
  wire [2:0] mem_0_1_mc;
  wire [1:0] mem_0_1_wa;
  wire [1:0] mem_0_1_wpulse;
  wire  mem_0_1_wpulseen;
  wire  mem_0_1_fwen;
  wire  mem_0_1_clkbyp;
  wire [8:0] mem_0_2_adr;
  wire  mem_0_2_clk;
  wire [63:0] mem_0_2_din;
  wire [63:0] mem_0_2_q;
  wire  mem_0_2_ren;
  wire  mem_0_2_wen;
  wire [63:0] mem_0_2_wbeb;
  wire  mem_0_2_mcen;
  wire [2:0] mem_0_2_mc;
  wire [1:0] mem_0_2_wa;
  wire [1:0] mem_0_2_wpulse;
  wire  mem_0_2_wpulseen;
  wire  mem_0_2_fwen;
  wire  mem_0_2_clkbyp;
  wire [8:0] mem_0_3_adr;
  wire  mem_0_3_clk;
  wire [63:0] mem_0_3_din;
  wire [63:0] mem_0_3_q;
  wire  mem_0_3_ren;
  wire  mem_0_3_wen;
  wire [63:0] mem_0_3_wbeb;
  wire  mem_0_3_mcen;
  wire [2:0] mem_0_3_mc;
  wire [1:0] mem_0_3_wa;
  wire [1:0] mem_0_3_wpulse;
  wire  mem_0_3_wpulseen;
  wire  mem_0_3_fwen;
  wire  mem_0_3_clkbyp;
  wire [63:0] RW0_rdata_0_0 = mem_0_0_q;
  wire [63:0] RW0_rdata_0_1 = mem_0_1_q;
  wire [63:0] RW0_rdata_0_2 = mem_0_2_q;
  wire [63:0] RW0_rdata_0_3 = mem_0_3_q;
  wire [127:0] _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [191:0] _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [255:0] RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire [127:0] _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire [191:0] _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0};
  wire  _GEN_4 = ~RW0_wmode;
  wire  _GEN_5 = RW0_wmask[0];
  wire  _GEN_6 = RW0_wmask[0];
  wire  _GEN_7 = RW0_wmask[0];
  wire [1:0] _GEN_8 = {RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_9 = RW0_wmask[0];
  wire [2:0] _GEN_10 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_11 = RW0_wmask[0];
  wire [3:0] _GEN_12 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_13 = RW0_wmask[0];
  wire [4:0] _GEN_14 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_15 = RW0_wmask[0];
  wire [5:0] _GEN_16 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_17 = RW0_wmask[0];
  wire [6:0] _GEN_18 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_19 = RW0_wmask[1];
  wire [7:0] _GEN_20 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0]};
  wire  _GEN_21 = RW0_wmask[1];
  wire [8:0] _GEN_22 = {RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_23 = RW0_wmask[1];
  wire [9:0] _GEN_24 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_25 = RW0_wmask[1];
  wire [10:0] _GEN_26 = {RW0_wmask[1],_GEN_24};
  wire  _GEN_27 = RW0_wmask[1];
  wire [11:0] _GEN_28 = {RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_29 = RW0_wmask[1];
  wire [12:0] _GEN_30 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_31 = RW0_wmask[1];
  wire [13:0] _GEN_32 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_33 = RW0_wmask[1];
  wire [14:0] _GEN_34 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_35 = RW0_wmask[2];
  wire [15:0] _GEN_36 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_37 = RW0_wmask[2];
  wire [16:0] _GEN_38 = {RW0_wmask[2],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    _GEN_24};
  wire  _GEN_39 = RW0_wmask[2];
  wire [17:0] _GEN_40 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],_GEN_24};
  wire  _GEN_41 = RW0_wmask[2];
  wire [18:0] _GEN_42 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],RW0_wmask[1],_GEN_24};
  wire  _GEN_43 = RW0_wmask[2];
  wire [19:0] _GEN_44 = {RW0_wmask[2],_GEN_42};
  wire  _GEN_45 = RW0_wmask[2];
  wire [20:0] _GEN_46 = {RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_47 = RW0_wmask[2];
  wire [21:0] _GEN_48 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_49 = RW0_wmask[2];
  wire [22:0] _GEN_50 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_51 = RW0_wmask[3];
  wire [23:0] _GEN_52 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_53 = RW0_wmask[3];
  wire [24:0] _GEN_54 = {RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_55 = RW0_wmask[3];
  wire [25:0] _GEN_56 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    _GEN_42};
  wire  _GEN_57 = RW0_wmask[3];
  wire [26:0] _GEN_58 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],_GEN_42};
  wire  _GEN_59 = RW0_wmask[3];
  wire [27:0] _GEN_60 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],RW0_wmask[2],_GEN_42};
  wire  _GEN_61 = RW0_wmask[3];
  wire [28:0] _GEN_62 = {RW0_wmask[3],_GEN_60};
  wire  _GEN_63 = RW0_wmask[3];
  wire [29:0] _GEN_64 = {RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_65 = RW0_wmask[3];
  wire [30:0] _GEN_66 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_67 = RW0_wmask[4];
  wire [31:0] _GEN_68 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_69 = RW0_wmask[4];
  wire [32:0] _GEN_70 = {RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_71 = RW0_wmask[4];
  wire [33:0] _GEN_72 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_73 = RW0_wmask[4];
  wire [34:0] _GEN_74 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    _GEN_60};
  wire  _GEN_75 = RW0_wmask[4];
  wire [35:0] _GEN_76 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],_GEN_60};
  wire  _GEN_77 = RW0_wmask[4];
  wire [36:0] _GEN_78 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],RW0_wmask[3],_GEN_60};
  wire  _GEN_79 = RW0_wmask[4];
  wire [37:0] _GEN_80 = {RW0_wmask[4],_GEN_78};
  wire  _GEN_81 = RW0_wmask[4];
  wire [38:0] _GEN_82 = {RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_83 = RW0_wmask[5];
  wire [39:0] _GEN_84 = {RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_85 = RW0_wmask[5];
  wire [40:0] _GEN_86 = {RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_87 = RW0_wmask[5];
  wire [41:0] _GEN_88 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_89 = RW0_wmask[5];
  wire [42:0] _GEN_90 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_91 = RW0_wmask[5];
  wire [43:0] _GEN_92 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],RW0_wmask[4],
    _GEN_78};
  wire  _GEN_93 = RW0_wmask[5];
  wire [44:0] _GEN_94 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],RW0_wmask[4],
    RW0_wmask[4],_GEN_78};
  wire  _GEN_95 = RW0_wmask[5];
  wire [45:0] _GEN_96 = {RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[5],RW0_wmask[4],
    RW0_wmask[4],RW0_wmask[4],_GEN_78};
  wire  _GEN_97 = RW0_wmask[5];
  wire [46:0] _GEN_98 = {RW0_wmask[5],_GEN_96};
  wire  _GEN_99 = RW0_wmask[6];
  wire [47:0] _GEN_100 = {RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_101 = RW0_wmask[6];
  wire [48:0] _GEN_102 = {RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_103 = RW0_wmask[6];
  wire [49:0] _GEN_104 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_105 = RW0_wmask[6];
  wire [50:0] _GEN_106 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_107 = RW0_wmask[6];
  wire [51:0] _GEN_108 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_109 = RW0_wmask[6];
  wire [52:0] _GEN_110 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],RW0_wmask[5],
    _GEN_96};
  wire  _GEN_111 = RW0_wmask[6];
  wire [53:0] _GEN_112 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[5],
    RW0_wmask[5],_GEN_96};
  wire  _GEN_113 = RW0_wmask[6];
  wire [54:0] _GEN_114 = {RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],RW0_wmask[6],
    RW0_wmask[5],RW0_wmask[5],_GEN_96};
  wire  _GEN_115 = RW0_wmask[7];
  wire [55:0] _GEN_116 = {RW0_wmask[6],_GEN_114};
  wire  _GEN_117 = RW0_wmask[7];
  wire [56:0] _GEN_118 = {RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_119 = RW0_wmask[7];
  wire [57:0] _GEN_120 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_121 = RW0_wmask[7];
  wire [58:0] _GEN_122 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_123 = RW0_wmask[7];
  wire [59:0] _GEN_124 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_125 = RW0_wmask[7];
  wire [60:0] _GEN_126 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_127 = RW0_wmask[7];
  wire [61:0] _GEN_128 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[6],
    _GEN_114};
  wire  _GEN_129 = RW0_wmask[7];
  wire [62:0] _GEN_130 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],
    RW0_wmask[6],_GEN_114};
  wire [63:0] _GEN_131 = {RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],RW0_wmask[7],
    RW0_wmask[7],RW0_wmask[6],_GEN_114};
  wire  _GEN_132 = ~RW0_wmode;
  wire  _GEN_133 = RW0_wmask[8];
  wire  _GEN_134 = RW0_wmask[8];
  wire  _GEN_135 = RW0_wmask[8];
  wire [1:0] _GEN_136 = {RW0_wmask[8],RW0_wmask[8]};
  wire  _GEN_137 = RW0_wmask[8];
  wire [2:0] _GEN_138 = {RW0_wmask[8],RW0_wmask[8],RW0_wmask[8]};
  wire  _GEN_139 = RW0_wmask[8];
  wire [3:0] _GEN_140 = {RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8]};
  wire  _GEN_141 = RW0_wmask[8];
  wire [4:0] _GEN_142 = {RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8]};
  wire  _GEN_143 = RW0_wmask[8];
  wire [5:0] _GEN_144 = {RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8]};
  wire  _GEN_145 = RW0_wmask[8];
  wire [6:0] _GEN_146 = {RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8]};
  wire  _GEN_147 = RW0_wmask[9];
  wire [7:0] _GEN_148 = {RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],
    RW0_wmask[8]};
  wire  _GEN_149 = RW0_wmask[9];
  wire [8:0] _GEN_150 = {RW0_wmask[9],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],
    RW0_wmask[8],RW0_wmask[8]};
  wire  _GEN_151 = RW0_wmask[9];
  wire [9:0] _GEN_152 = {RW0_wmask[9],RW0_wmask[9],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],RW0_wmask[8],
    RW0_wmask[8],RW0_wmask[8],RW0_wmask[8]};
  wire  _GEN_153 = RW0_wmask[9];
  wire [10:0] _GEN_154 = {RW0_wmask[9],_GEN_152};
  wire  _GEN_155 = RW0_wmask[9];
  wire [11:0] _GEN_156 = {RW0_wmask[9],RW0_wmask[9],_GEN_152};
  wire  _GEN_157 = RW0_wmask[9];
  wire [12:0] _GEN_158 = {RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],_GEN_152};
  wire  _GEN_159 = RW0_wmask[9];
  wire [13:0] _GEN_160 = {RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],_GEN_152};
  wire  _GEN_161 = RW0_wmask[9];
  wire [14:0] _GEN_162 = {RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],_GEN_152};
  wire  _GEN_163 = RW0_wmask[10];
  wire [15:0] _GEN_164 = {RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],_GEN_152};
  wire  _GEN_165 = RW0_wmask[10];
  wire [16:0] _GEN_166 = {RW0_wmask[10],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],
    _GEN_152};
  wire  _GEN_167 = RW0_wmask[10];
  wire [17:0] _GEN_168 = {RW0_wmask[10],RW0_wmask[10],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],
    RW0_wmask[9],_GEN_152};
  wire  _GEN_169 = RW0_wmask[10];
  wire [18:0] _GEN_170 = {RW0_wmask[10],RW0_wmask[10],RW0_wmask[10],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],RW0_wmask[9],
    RW0_wmask[9],RW0_wmask[9],_GEN_152};
  wire  _GEN_171 = RW0_wmask[10];
  wire [19:0] _GEN_172 = {RW0_wmask[10],_GEN_170};
  wire  _GEN_173 = RW0_wmask[10];
  wire [20:0] _GEN_174 = {RW0_wmask[10],RW0_wmask[10],_GEN_170};
  wire  _GEN_175 = RW0_wmask[10];
  wire [21:0] _GEN_176 = {RW0_wmask[10],RW0_wmask[10],RW0_wmask[10],_GEN_170};
  wire  _GEN_177 = RW0_wmask[10];
  wire [22:0] _GEN_178 = {RW0_wmask[10],RW0_wmask[10],RW0_wmask[10],RW0_wmask[10],_GEN_170};
  wire  _GEN_179 = RW0_wmask[11];
  wire [23:0] _GEN_180 = {RW0_wmask[10],RW0_wmask[10],RW0_wmask[10],RW0_wmask[10],RW0_wmask[10],_GEN_170};
  wire  _GEN_181 = RW0_wmask[11];
  wire [24:0] _GEN_182 = {RW0_wmask[11],RW0_wmask[10],RW0_wmask[10],RW0_wmask[10],RW0_wmask[10],RW0_wmask[10],_GEN_170};
  wire  _GEN_183 = RW0_wmask[11];
  wire [25:0] _GEN_184 = {RW0_wmask[11],RW0_wmask[11],RW0_wmask[10],RW0_wmask[10],RW0_wmask[10],RW0_wmask[10],RW0_wmask[
    10],_GEN_170};
  wire  _GEN_185 = RW0_wmask[11];
  wire [26:0] _GEN_186 = {RW0_wmask[11],RW0_wmask[11],RW0_wmask[11],RW0_wmask[10],RW0_wmask[10],RW0_wmask[10],RW0_wmask[
    10],RW0_wmask[10],_GEN_170};
  wire  _GEN_187 = RW0_wmask[11];
  wire [27:0] _GEN_188 = {RW0_wmask[11],RW0_wmask[11],RW0_wmask[11],RW0_wmask[11],RW0_wmask[10],RW0_wmask[10],RW0_wmask[
    10],RW0_wmask[10],RW0_wmask[10],_GEN_170};
  wire  _GEN_189 = RW0_wmask[11];
  wire [28:0] _GEN_190 = {RW0_wmask[11],_GEN_188};
  wire  _GEN_191 = RW0_wmask[11];
  wire [29:0] _GEN_192 = {RW0_wmask[11],RW0_wmask[11],_GEN_188};
  wire  _GEN_193 = RW0_wmask[11];
  wire [30:0] _GEN_194 = {RW0_wmask[11],RW0_wmask[11],RW0_wmask[11],_GEN_188};
  wire  _GEN_195 = RW0_wmask[12];
  wire [31:0] _GEN_196 = {RW0_wmask[11],RW0_wmask[11],RW0_wmask[11],RW0_wmask[11],_GEN_188};
  wire  _GEN_197 = RW0_wmask[12];
  wire [32:0] _GEN_198 = {RW0_wmask[12],RW0_wmask[11],RW0_wmask[11],RW0_wmask[11],RW0_wmask[11],_GEN_188};
  wire  _GEN_199 = RW0_wmask[12];
  wire [33:0] _GEN_200 = {RW0_wmask[12],RW0_wmask[12],RW0_wmask[11],RW0_wmask[11],RW0_wmask[11],RW0_wmask[11],_GEN_188};
  wire  _GEN_201 = RW0_wmask[12];
  wire [34:0] _GEN_202 = {RW0_wmask[12],RW0_wmask[12],RW0_wmask[12],RW0_wmask[11],RW0_wmask[11],RW0_wmask[11],RW0_wmask[
    11],_GEN_188};
  wire  _GEN_203 = RW0_wmask[12];
  wire [35:0] _GEN_204 = {RW0_wmask[12],RW0_wmask[12],RW0_wmask[12],RW0_wmask[12],RW0_wmask[11],RW0_wmask[11],RW0_wmask[
    11],RW0_wmask[11],_GEN_188};
  wire  _GEN_205 = RW0_wmask[12];
  wire [36:0] _GEN_206 = {RW0_wmask[12],RW0_wmask[12],RW0_wmask[12],RW0_wmask[12],RW0_wmask[12],RW0_wmask[11],RW0_wmask[
    11],RW0_wmask[11],RW0_wmask[11],_GEN_188};
  wire  _GEN_207 = RW0_wmask[12];
  wire [37:0] _GEN_208 = {RW0_wmask[12],_GEN_206};
  wire  _GEN_209 = RW0_wmask[12];
  wire [38:0] _GEN_210 = {RW0_wmask[12],RW0_wmask[12],_GEN_206};
  wire  _GEN_211 = RW0_wmask[13];
  wire [39:0] _GEN_212 = {RW0_wmask[12],RW0_wmask[12],RW0_wmask[12],_GEN_206};
  wire  _GEN_213 = RW0_wmask[13];
  wire [40:0] _GEN_214 = {RW0_wmask[13],RW0_wmask[12],RW0_wmask[12],RW0_wmask[12],_GEN_206};
  wire  _GEN_215 = RW0_wmask[13];
  wire [41:0] _GEN_216 = {RW0_wmask[13],RW0_wmask[13],RW0_wmask[12],RW0_wmask[12],RW0_wmask[12],_GEN_206};
  wire  _GEN_217 = RW0_wmask[13];
  wire [42:0] _GEN_218 = {RW0_wmask[13],RW0_wmask[13],RW0_wmask[13],RW0_wmask[12],RW0_wmask[12],RW0_wmask[12],_GEN_206};
  wire  _GEN_219 = RW0_wmask[13];
  wire [43:0] _GEN_220 = {RW0_wmask[13],RW0_wmask[13],RW0_wmask[13],RW0_wmask[13],RW0_wmask[12],RW0_wmask[12],RW0_wmask[
    12],_GEN_206};
  wire  _GEN_221 = RW0_wmask[13];
  wire [44:0] _GEN_222 = {RW0_wmask[13],RW0_wmask[13],RW0_wmask[13],RW0_wmask[13],RW0_wmask[13],RW0_wmask[12],RW0_wmask[
    12],RW0_wmask[12],_GEN_206};
  wire  _GEN_223 = RW0_wmask[13];
  wire [45:0] _GEN_224 = {RW0_wmask[13],RW0_wmask[13],RW0_wmask[13],RW0_wmask[13],RW0_wmask[13],RW0_wmask[13],RW0_wmask[
    12],RW0_wmask[12],RW0_wmask[12],_GEN_206};
  wire  _GEN_225 = RW0_wmask[13];
  wire [46:0] _GEN_226 = {RW0_wmask[13],_GEN_224};
  wire  _GEN_227 = RW0_wmask[14];
  wire [47:0] _GEN_228 = {RW0_wmask[13],RW0_wmask[13],_GEN_224};
  wire  _GEN_229 = RW0_wmask[14];
  wire [48:0] _GEN_230 = {RW0_wmask[14],RW0_wmask[13],RW0_wmask[13],_GEN_224};
  wire  _GEN_231 = RW0_wmask[14];
  wire [49:0] _GEN_232 = {RW0_wmask[14],RW0_wmask[14],RW0_wmask[13],RW0_wmask[13],_GEN_224};
  wire  _GEN_233 = RW0_wmask[14];
  wire [50:0] _GEN_234 = {RW0_wmask[14],RW0_wmask[14],RW0_wmask[14],RW0_wmask[13],RW0_wmask[13],_GEN_224};
  wire  _GEN_235 = RW0_wmask[14];
  wire [51:0] _GEN_236 = {RW0_wmask[14],RW0_wmask[14],RW0_wmask[14],RW0_wmask[14],RW0_wmask[13],RW0_wmask[13],_GEN_224};
  wire  _GEN_237 = RW0_wmask[14];
  wire [52:0] _GEN_238 = {RW0_wmask[14],RW0_wmask[14],RW0_wmask[14],RW0_wmask[14],RW0_wmask[14],RW0_wmask[13],RW0_wmask[
    13],_GEN_224};
  wire  _GEN_239 = RW0_wmask[14];
  wire [53:0] _GEN_240 = {RW0_wmask[14],RW0_wmask[14],RW0_wmask[14],RW0_wmask[14],RW0_wmask[14],RW0_wmask[14],RW0_wmask[
    13],RW0_wmask[13],_GEN_224};
  wire  _GEN_241 = RW0_wmask[14];
  wire [54:0] _GEN_242 = {RW0_wmask[14],RW0_wmask[14],RW0_wmask[14],RW0_wmask[14],RW0_wmask[14],RW0_wmask[14],RW0_wmask[
    14],RW0_wmask[13],RW0_wmask[13],_GEN_224};
  wire  _GEN_243 = RW0_wmask[15];
  wire [55:0] _GEN_244 = {RW0_wmask[14],_GEN_242};
  wire  _GEN_245 = RW0_wmask[15];
  wire [56:0] _GEN_246 = {RW0_wmask[15],RW0_wmask[14],_GEN_242};
  wire  _GEN_247 = RW0_wmask[15];
  wire [57:0] _GEN_248 = {RW0_wmask[15],RW0_wmask[15],RW0_wmask[14],_GEN_242};
  wire  _GEN_249 = RW0_wmask[15];
  wire [58:0] _GEN_250 = {RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[14],_GEN_242};
  wire  _GEN_251 = RW0_wmask[15];
  wire [59:0] _GEN_252 = {RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[14],_GEN_242};
  wire  _GEN_253 = RW0_wmask[15];
  wire [60:0] _GEN_254 = {RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[14],_GEN_242};
  wire  _GEN_255 = RW0_wmask[15];
  wire [61:0] _GEN_256 = {RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[
    14],_GEN_242};
  wire  _GEN_257 = RW0_wmask[15];
  wire [62:0] _GEN_258 = {RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[
    15],RW0_wmask[14],_GEN_242};
  wire [63:0] _GEN_259 = {RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[15],RW0_wmask[
    15],RW0_wmask[15],RW0_wmask[14],_GEN_242};
  wire  _GEN_260 = ~RW0_wmode;
  wire  _GEN_261 = RW0_wmask[16];
  wire  _GEN_262 = RW0_wmask[16];
  wire  _GEN_263 = RW0_wmask[16];
  wire [1:0] _GEN_264 = {RW0_wmask[16],RW0_wmask[16]};
  wire  _GEN_265 = RW0_wmask[16];
  wire [2:0] _GEN_266 = {RW0_wmask[16],RW0_wmask[16],RW0_wmask[16]};
  wire  _GEN_267 = RW0_wmask[16];
  wire [3:0] _GEN_268 = {RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16]};
  wire  _GEN_269 = RW0_wmask[16];
  wire [4:0] _GEN_270 = {RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16]};
  wire  _GEN_271 = RW0_wmask[16];
  wire [5:0] _GEN_272 = {RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16]};
  wire  _GEN_273 = RW0_wmask[16];
  wire [6:0] _GEN_274 = {RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[
    16]};
  wire  _GEN_275 = RW0_wmask[17];
  wire [7:0] _GEN_276 = {RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[
    16],RW0_wmask[16]};
  wire  _GEN_277 = RW0_wmask[17];
  wire [8:0] _GEN_278 = {RW0_wmask[17],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[
    16],RW0_wmask[16],RW0_wmask[16]};
  wire  _GEN_279 = RW0_wmask[17];
  wire [9:0] _GEN_280 = {RW0_wmask[17],RW0_wmask[17],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[
    16],RW0_wmask[16],RW0_wmask[16],RW0_wmask[16]};
  wire  _GEN_281 = RW0_wmask[17];
  wire [10:0] _GEN_282 = {RW0_wmask[17],_GEN_280};
  wire  _GEN_283 = RW0_wmask[17];
  wire [11:0] _GEN_284 = {RW0_wmask[17],RW0_wmask[17],_GEN_280};
  wire  _GEN_285 = RW0_wmask[17];
  wire [12:0] _GEN_286 = {RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],_GEN_280};
  wire  _GEN_287 = RW0_wmask[17];
  wire [13:0] _GEN_288 = {RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],_GEN_280};
  wire  _GEN_289 = RW0_wmask[17];
  wire [14:0] _GEN_290 = {RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],_GEN_280};
  wire  _GEN_291 = RW0_wmask[18];
  wire [15:0] _GEN_292 = {RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],_GEN_280};
  wire  _GEN_293 = RW0_wmask[18];
  wire [16:0] _GEN_294 = {RW0_wmask[18],RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],RW0_wmask[
    17],_GEN_280};
  wire  _GEN_295 = RW0_wmask[18];
  wire [17:0] _GEN_296 = {RW0_wmask[18],RW0_wmask[18],RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],RW0_wmask[
    17],RW0_wmask[17],_GEN_280};
  wire  _GEN_297 = RW0_wmask[18];
  wire [18:0] _GEN_298 = {RW0_wmask[18],RW0_wmask[18],RW0_wmask[18],RW0_wmask[17],RW0_wmask[17],RW0_wmask[17],RW0_wmask[
    17],RW0_wmask[17],RW0_wmask[17],_GEN_280};
  wire  _GEN_299 = RW0_wmask[18];
  wire [19:0] _GEN_300 = {RW0_wmask[18],_GEN_298};
  wire  _GEN_301 = RW0_wmask[18];
  wire [20:0] _GEN_302 = {RW0_wmask[18],RW0_wmask[18],_GEN_298};
  wire  _GEN_303 = RW0_wmask[18];
  wire [21:0] _GEN_304 = {RW0_wmask[18],RW0_wmask[18],RW0_wmask[18],_GEN_298};
  wire  _GEN_305 = RW0_wmask[18];
  wire [22:0] _GEN_306 = {RW0_wmask[18],RW0_wmask[18],RW0_wmask[18],RW0_wmask[18],_GEN_298};
  wire  _GEN_307 = RW0_wmask[19];
  wire [23:0] _GEN_308 = {RW0_wmask[18],RW0_wmask[18],RW0_wmask[18],RW0_wmask[18],RW0_wmask[18],_GEN_298};
  wire  _GEN_309 = RW0_wmask[19];
  wire [24:0] _GEN_310 = {RW0_wmask[19],RW0_wmask[18],RW0_wmask[18],RW0_wmask[18],RW0_wmask[18],RW0_wmask[18],_GEN_298};
  wire  _GEN_311 = RW0_wmask[19];
  wire [25:0] _GEN_312 = {RW0_wmask[19],RW0_wmask[19],RW0_wmask[18],RW0_wmask[18],RW0_wmask[18],RW0_wmask[18],RW0_wmask[
    18],_GEN_298};
  wire  _GEN_313 = RW0_wmask[19];
  wire [26:0] _GEN_314 = {RW0_wmask[19],RW0_wmask[19],RW0_wmask[19],RW0_wmask[18],RW0_wmask[18],RW0_wmask[18],RW0_wmask[
    18],RW0_wmask[18],_GEN_298};
  wire  _GEN_315 = RW0_wmask[19];
  wire [27:0] _GEN_316 = {RW0_wmask[19],RW0_wmask[19],RW0_wmask[19],RW0_wmask[19],RW0_wmask[18],RW0_wmask[18],RW0_wmask[
    18],RW0_wmask[18],RW0_wmask[18],_GEN_298};
  wire  _GEN_317 = RW0_wmask[19];
  wire [28:0] _GEN_318 = {RW0_wmask[19],_GEN_316};
  wire  _GEN_319 = RW0_wmask[19];
  wire [29:0] _GEN_320 = {RW0_wmask[19],RW0_wmask[19],_GEN_316};
  wire  _GEN_321 = RW0_wmask[19];
  wire [30:0] _GEN_322 = {RW0_wmask[19],RW0_wmask[19],RW0_wmask[19],_GEN_316};
  wire  _GEN_323 = RW0_wmask[20];
  wire [31:0] _GEN_324 = {RW0_wmask[19],RW0_wmask[19],RW0_wmask[19],RW0_wmask[19],_GEN_316};
  wire  _GEN_325 = RW0_wmask[20];
  wire [32:0] _GEN_326 = {RW0_wmask[20],RW0_wmask[19],RW0_wmask[19],RW0_wmask[19],RW0_wmask[19],_GEN_316};
  wire  _GEN_327 = RW0_wmask[20];
  wire [33:0] _GEN_328 = {RW0_wmask[20],RW0_wmask[20],RW0_wmask[19],RW0_wmask[19],RW0_wmask[19],RW0_wmask[19],_GEN_316};
  wire  _GEN_329 = RW0_wmask[20];
  wire [34:0] _GEN_330 = {RW0_wmask[20],RW0_wmask[20],RW0_wmask[20],RW0_wmask[19],RW0_wmask[19],RW0_wmask[19],RW0_wmask[
    19],_GEN_316};
  wire  _GEN_331 = RW0_wmask[20];
  wire [35:0] _GEN_332 = {RW0_wmask[20],RW0_wmask[20],RW0_wmask[20],RW0_wmask[20],RW0_wmask[19],RW0_wmask[19],RW0_wmask[
    19],RW0_wmask[19],_GEN_316};
  wire  _GEN_333 = RW0_wmask[20];
  wire [36:0] _GEN_334 = {RW0_wmask[20],RW0_wmask[20],RW0_wmask[20],RW0_wmask[20],RW0_wmask[20],RW0_wmask[19],RW0_wmask[
    19],RW0_wmask[19],RW0_wmask[19],_GEN_316};
  wire  _GEN_335 = RW0_wmask[20];
  wire [37:0] _GEN_336 = {RW0_wmask[20],_GEN_334};
  wire  _GEN_337 = RW0_wmask[20];
  wire [38:0] _GEN_338 = {RW0_wmask[20],RW0_wmask[20],_GEN_334};
  wire  _GEN_339 = RW0_wmask[21];
  wire [39:0] _GEN_340 = {RW0_wmask[20],RW0_wmask[20],RW0_wmask[20],_GEN_334};
  wire  _GEN_341 = RW0_wmask[21];
  wire [40:0] _GEN_342 = {RW0_wmask[21],RW0_wmask[20],RW0_wmask[20],RW0_wmask[20],_GEN_334};
  wire  _GEN_343 = RW0_wmask[21];
  wire [41:0] _GEN_344 = {RW0_wmask[21],RW0_wmask[21],RW0_wmask[20],RW0_wmask[20],RW0_wmask[20],_GEN_334};
  wire  _GEN_345 = RW0_wmask[21];
  wire [42:0] _GEN_346 = {RW0_wmask[21],RW0_wmask[21],RW0_wmask[21],RW0_wmask[20],RW0_wmask[20],RW0_wmask[20],_GEN_334};
  wire  _GEN_347 = RW0_wmask[21];
  wire [43:0] _GEN_348 = {RW0_wmask[21],RW0_wmask[21],RW0_wmask[21],RW0_wmask[21],RW0_wmask[20],RW0_wmask[20],RW0_wmask[
    20],_GEN_334};
  wire  _GEN_349 = RW0_wmask[21];
  wire [44:0] _GEN_350 = {RW0_wmask[21],RW0_wmask[21],RW0_wmask[21],RW0_wmask[21],RW0_wmask[21],RW0_wmask[20],RW0_wmask[
    20],RW0_wmask[20],_GEN_334};
  wire  _GEN_351 = RW0_wmask[21];
  wire [45:0] _GEN_352 = {RW0_wmask[21],RW0_wmask[21],RW0_wmask[21],RW0_wmask[21],RW0_wmask[21],RW0_wmask[21],RW0_wmask[
    20],RW0_wmask[20],RW0_wmask[20],_GEN_334};
  wire  _GEN_353 = RW0_wmask[21];
  wire [46:0] _GEN_354 = {RW0_wmask[21],_GEN_352};
  wire  _GEN_355 = RW0_wmask[22];
  wire [47:0] _GEN_356 = {RW0_wmask[21],RW0_wmask[21],_GEN_352};
  wire  _GEN_357 = RW0_wmask[22];
  wire [48:0] _GEN_358 = {RW0_wmask[22],RW0_wmask[21],RW0_wmask[21],_GEN_352};
  wire  _GEN_359 = RW0_wmask[22];
  wire [49:0] _GEN_360 = {RW0_wmask[22],RW0_wmask[22],RW0_wmask[21],RW0_wmask[21],_GEN_352};
  wire  _GEN_361 = RW0_wmask[22];
  wire [50:0] _GEN_362 = {RW0_wmask[22],RW0_wmask[22],RW0_wmask[22],RW0_wmask[21],RW0_wmask[21],_GEN_352};
  wire  _GEN_363 = RW0_wmask[22];
  wire [51:0] _GEN_364 = {RW0_wmask[22],RW0_wmask[22],RW0_wmask[22],RW0_wmask[22],RW0_wmask[21],RW0_wmask[21],_GEN_352};
  wire  _GEN_365 = RW0_wmask[22];
  wire [52:0] _GEN_366 = {RW0_wmask[22],RW0_wmask[22],RW0_wmask[22],RW0_wmask[22],RW0_wmask[22],RW0_wmask[21],RW0_wmask[
    21],_GEN_352};
  wire  _GEN_367 = RW0_wmask[22];
  wire [53:0] _GEN_368 = {RW0_wmask[22],RW0_wmask[22],RW0_wmask[22],RW0_wmask[22],RW0_wmask[22],RW0_wmask[22],RW0_wmask[
    21],RW0_wmask[21],_GEN_352};
  wire  _GEN_369 = RW0_wmask[22];
  wire [54:0] _GEN_370 = {RW0_wmask[22],RW0_wmask[22],RW0_wmask[22],RW0_wmask[22],RW0_wmask[22],RW0_wmask[22],RW0_wmask[
    22],RW0_wmask[21],RW0_wmask[21],_GEN_352};
  wire  _GEN_371 = RW0_wmask[23];
  wire [55:0] _GEN_372 = {RW0_wmask[22],_GEN_370};
  wire  _GEN_373 = RW0_wmask[23];
  wire [56:0] _GEN_374 = {RW0_wmask[23],RW0_wmask[22],_GEN_370};
  wire  _GEN_375 = RW0_wmask[23];
  wire [57:0] _GEN_376 = {RW0_wmask[23],RW0_wmask[23],RW0_wmask[22],_GEN_370};
  wire  _GEN_377 = RW0_wmask[23];
  wire [58:0] _GEN_378 = {RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[22],_GEN_370};
  wire  _GEN_379 = RW0_wmask[23];
  wire [59:0] _GEN_380 = {RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[22],_GEN_370};
  wire  _GEN_381 = RW0_wmask[23];
  wire [60:0] _GEN_382 = {RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[22],_GEN_370};
  wire  _GEN_383 = RW0_wmask[23];
  wire [61:0] _GEN_384 = {RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[
    22],_GEN_370};
  wire  _GEN_385 = RW0_wmask[23];
  wire [62:0] _GEN_386 = {RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[
    23],RW0_wmask[22],_GEN_370};
  wire [63:0] _GEN_387 = {RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[23],RW0_wmask[
    23],RW0_wmask[23],RW0_wmask[22],_GEN_370};
  wire  _GEN_388 = ~RW0_wmode;
  wire  _GEN_389 = RW0_wmask[24];
  wire  _GEN_390 = RW0_wmask[24];
  wire  _GEN_391 = RW0_wmask[24];
  wire [1:0] _GEN_392 = {RW0_wmask[24],RW0_wmask[24]};
  wire  _GEN_393 = RW0_wmask[24];
  wire [2:0] _GEN_394 = {RW0_wmask[24],RW0_wmask[24],RW0_wmask[24]};
  wire  _GEN_395 = RW0_wmask[24];
  wire [3:0] _GEN_396 = {RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24]};
  wire  _GEN_397 = RW0_wmask[24];
  wire [4:0] _GEN_398 = {RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24]};
  wire  _GEN_399 = RW0_wmask[24];
  wire [5:0] _GEN_400 = {RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24]};
  wire  _GEN_401 = RW0_wmask[24];
  wire [6:0] _GEN_402 = {RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[
    24]};
  wire  _GEN_403 = RW0_wmask[25];
  wire [7:0] _GEN_404 = {RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[
    24],RW0_wmask[24]};
  wire  _GEN_405 = RW0_wmask[25];
  wire [8:0] _GEN_406 = {RW0_wmask[25],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[
    24],RW0_wmask[24],RW0_wmask[24]};
  wire  _GEN_407 = RW0_wmask[25];
  wire [9:0] _GEN_408 = {RW0_wmask[25],RW0_wmask[25],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[
    24],RW0_wmask[24],RW0_wmask[24],RW0_wmask[24]};
  wire  _GEN_409 = RW0_wmask[25];
  wire [10:0] _GEN_410 = {RW0_wmask[25],_GEN_408};
  wire  _GEN_411 = RW0_wmask[25];
  wire [11:0] _GEN_412 = {RW0_wmask[25],RW0_wmask[25],_GEN_408};
  wire  _GEN_413 = RW0_wmask[25];
  wire [12:0] _GEN_414 = {RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],_GEN_408};
  wire  _GEN_415 = RW0_wmask[25];
  wire [13:0] _GEN_416 = {RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],_GEN_408};
  wire  _GEN_417 = RW0_wmask[25];
  wire [14:0] _GEN_418 = {RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],_GEN_408};
  wire  _GEN_419 = RW0_wmask[26];
  wire [15:0] _GEN_420 = {RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],_GEN_408};
  wire  _GEN_421 = RW0_wmask[26];
  wire [16:0] _GEN_422 = {RW0_wmask[26],RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],RW0_wmask[
    25],_GEN_408};
  wire  _GEN_423 = RW0_wmask[26];
  wire [17:0] _GEN_424 = {RW0_wmask[26],RW0_wmask[26],RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],RW0_wmask[
    25],RW0_wmask[25],_GEN_408};
  wire  _GEN_425 = RW0_wmask[26];
  wire [18:0] _GEN_426 = {RW0_wmask[26],RW0_wmask[26],RW0_wmask[26],RW0_wmask[25],RW0_wmask[25],RW0_wmask[25],RW0_wmask[
    25],RW0_wmask[25],RW0_wmask[25],_GEN_408};
  wire  _GEN_427 = RW0_wmask[26];
  wire [19:0] _GEN_428 = {RW0_wmask[26],_GEN_426};
  wire  _GEN_429 = RW0_wmask[26];
  wire [20:0] _GEN_430 = {RW0_wmask[26],RW0_wmask[26],_GEN_426};
  wire  _GEN_431 = RW0_wmask[26];
  wire [21:0] _GEN_432 = {RW0_wmask[26],RW0_wmask[26],RW0_wmask[26],_GEN_426};
  wire  _GEN_433 = RW0_wmask[26];
  wire [22:0] _GEN_434 = {RW0_wmask[26],RW0_wmask[26],RW0_wmask[26],RW0_wmask[26],_GEN_426};
  wire  _GEN_435 = RW0_wmask[27];
  wire [23:0] _GEN_436 = {RW0_wmask[26],RW0_wmask[26],RW0_wmask[26],RW0_wmask[26],RW0_wmask[26],_GEN_426};
  wire  _GEN_437 = RW0_wmask[27];
  wire [24:0] _GEN_438 = {RW0_wmask[27],RW0_wmask[26],RW0_wmask[26],RW0_wmask[26],RW0_wmask[26],RW0_wmask[26],_GEN_426};
  wire  _GEN_439 = RW0_wmask[27];
  wire [25:0] _GEN_440 = {RW0_wmask[27],RW0_wmask[27],RW0_wmask[26],RW0_wmask[26],RW0_wmask[26],RW0_wmask[26],RW0_wmask[
    26],_GEN_426};
  wire  _GEN_441 = RW0_wmask[27];
  wire [26:0] _GEN_442 = {RW0_wmask[27],RW0_wmask[27],RW0_wmask[27],RW0_wmask[26],RW0_wmask[26],RW0_wmask[26],RW0_wmask[
    26],RW0_wmask[26],_GEN_426};
  wire  _GEN_443 = RW0_wmask[27];
  wire [27:0] _GEN_444 = {RW0_wmask[27],RW0_wmask[27],RW0_wmask[27],RW0_wmask[27],RW0_wmask[26],RW0_wmask[26],RW0_wmask[
    26],RW0_wmask[26],RW0_wmask[26],_GEN_426};
  wire  _GEN_445 = RW0_wmask[27];
  wire [28:0] _GEN_446 = {RW0_wmask[27],_GEN_444};
  wire  _GEN_447 = RW0_wmask[27];
  wire [29:0] _GEN_448 = {RW0_wmask[27],RW0_wmask[27],_GEN_444};
  wire  _GEN_449 = RW0_wmask[27];
  wire [30:0] _GEN_450 = {RW0_wmask[27],RW0_wmask[27],RW0_wmask[27],_GEN_444};
  wire  _GEN_451 = RW0_wmask[28];
  wire [31:0] _GEN_452 = {RW0_wmask[27],RW0_wmask[27],RW0_wmask[27],RW0_wmask[27],_GEN_444};
  wire  _GEN_453 = RW0_wmask[28];
  wire [32:0] _GEN_454 = {RW0_wmask[28],RW0_wmask[27],RW0_wmask[27],RW0_wmask[27],RW0_wmask[27],_GEN_444};
  wire  _GEN_455 = RW0_wmask[28];
  wire [33:0] _GEN_456 = {RW0_wmask[28],RW0_wmask[28],RW0_wmask[27],RW0_wmask[27],RW0_wmask[27],RW0_wmask[27],_GEN_444};
  wire  _GEN_457 = RW0_wmask[28];
  wire [34:0] _GEN_458 = {RW0_wmask[28],RW0_wmask[28],RW0_wmask[28],RW0_wmask[27],RW0_wmask[27],RW0_wmask[27],RW0_wmask[
    27],_GEN_444};
  wire  _GEN_459 = RW0_wmask[28];
  wire [35:0] _GEN_460 = {RW0_wmask[28],RW0_wmask[28],RW0_wmask[28],RW0_wmask[28],RW0_wmask[27],RW0_wmask[27],RW0_wmask[
    27],RW0_wmask[27],_GEN_444};
  wire  _GEN_461 = RW0_wmask[28];
  wire [36:0] _GEN_462 = {RW0_wmask[28],RW0_wmask[28],RW0_wmask[28],RW0_wmask[28],RW0_wmask[28],RW0_wmask[27],RW0_wmask[
    27],RW0_wmask[27],RW0_wmask[27],_GEN_444};
  wire  _GEN_463 = RW0_wmask[28];
  wire [37:0] _GEN_464 = {RW0_wmask[28],_GEN_462};
  wire  _GEN_465 = RW0_wmask[28];
  wire [38:0] _GEN_466 = {RW0_wmask[28],RW0_wmask[28],_GEN_462};
  wire  _GEN_467 = RW0_wmask[29];
  wire [39:0] _GEN_468 = {RW0_wmask[28],RW0_wmask[28],RW0_wmask[28],_GEN_462};
  wire  _GEN_469 = RW0_wmask[29];
  wire [40:0] _GEN_470 = {RW0_wmask[29],RW0_wmask[28],RW0_wmask[28],RW0_wmask[28],_GEN_462};
  wire  _GEN_471 = RW0_wmask[29];
  wire [41:0] _GEN_472 = {RW0_wmask[29],RW0_wmask[29],RW0_wmask[28],RW0_wmask[28],RW0_wmask[28],_GEN_462};
  wire  _GEN_473 = RW0_wmask[29];
  wire [42:0] _GEN_474 = {RW0_wmask[29],RW0_wmask[29],RW0_wmask[29],RW0_wmask[28],RW0_wmask[28],RW0_wmask[28],_GEN_462};
  wire  _GEN_475 = RW0_wmask[29];
  wire [43:0] _GEN_476 = {RW0_wmask[29],RW0_wmask[29],RW0_wmask[29],RW0_wmask[29],RW0_wmask[28],RW0_wmask[28],RW0_wmask[
    28],_GEN_462};
  wire  _GEN_477 = RW0_wmask[29];
  wire [44:0] _GEN_478 = {RW0_wmask[29],RW0_wmask[29],RW0_wmask[29],RW0_wmask[29],RW0_wmask[29],RW0_wmask[28],RW0_wmask[
    28],RW0_wmask[28],_GEN_462};
  wire  _GEN_479 = RW0_wmask[29];
  wire [45:0] _GEN_480 = {RW0_wmask[29],RW0_wmask[29],RW0_wmask[29],RW0_wmask[29],RW0_wmask[29],RW0_wmask[29],RW0_wmask[
    28],RW0_wmask[28],RW0_wmask[28],_GEN_462};
  wire  _GEN_481 = RW0_wmask[29];
  wire [46:0] _GEN_482 = {RW0_wmask[29],_GEN_480};
  wire  _GEN_483 = RW0_wmask[30];
  wire [47:0] _GEN_484 = {RW0_wmask[29],RW0_wmask[29],_GEN_480};
  wire  _GEN_485 = RW0_wmask[30];
  wire [48:0] _GEN_486 = {RW0_wmask[30],RW0_wmask[29],RW0_wmask[29],_GEN_480};
  wire  _GEN_487 = RW0_wmask[30];
  wire [49:0] _GEN_488 = {RW0_wmask[30],RW0_wmask[30],RW0_wmask[29],RW0_wmask[29],_GEN_480};
  wire  _GEN_489 = RW0_wmask[30];
  wire [50:0] _GEN_490 = {RW0_wmask[30],RW0_wmask[30],RW0_wmask[30],RW0_wmask[29],RW0_wmask[29],_GEN_480};
  wire  _GEN_491 = RW0_wmask[30];
  wire [51:0] _GEN_492 = {RW0_wmask[30],RW0_wmask[30],RW0_wmask[30],RW0_wmask[30],RW0_wmask[29],RW0_wmask[29],_GEN_480};
  wire  _GEN_493 = RW0_wmask[30];
  wire [52:0] _GEN_494 = {RW0_wmask[30],RW0_wmask[30],RW0_wmask[30],RW0_wmask[30],RW0_wmask[30],RW0_wmask[29],RW0_wmask[
    29],_GEN_480};
  wire  _GEN_495 = RW0_wmask[30];
  wire [53:0] _GEN_496 = {RW0_wmask[30],RW0_wmask[30],RW0_wmask[30],RW0_wmask[30],RW0_wmask[30],RW0_wmask[30],RW0_wmask[
    29],RW0_wmask[29],_GEN_480};
  wire  _GEN_497 = RW0_wmask[30];
  wire [54:0] _GEN_498 = {RW0_wmask[30],RW0_wmask[30],RW0_wmask[30],RW0_wmask[30],RW0_wmask[30],RW0_wmask[30],RW0_wmask[
    30],RW0_wmask[29],RW0_wmask[29],_GEN_480};
  wire  _GEN_499 = RW0_wmask[31];
  wire [55:0] _GEN_500 = {RW0_wmask[30],_GEN_498};
  wire  _GEN_501 = RW0_wmask[31];
  wire [56:0] _GEN_502 = {RW0_wmask[31],RW0_wmask[30],_GEN_498};
  wire  _GEN_503 = RW0_wmask[31];
  wire [57:0] _GEN_504 = {RW0_wmask[31],RW0_wmask[31],RW0_wmask[30],_GEN_498};
  wire  _GEN_505 = RW0_wmask[31];
  wire [58:0] _GEN_506 = {RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[30],_GEN_498};
  wire  _GEN_507 = RW0_wmask[31];
  wire [59:0] _GEN_508 = {RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[30],_GEN_498};
  wire  _GEN_509 = RW0_wmask[31];
  wire [60:0] _GEN_510 = {RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[30],_GEN_498};
  wire  _GEN_511 = RW0_wmask[31];
  wire [61:0] _GEN_512 = {RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[
    30],_GEN_498};
  wire  _GEN_513 = RW0_wmask[31];
  wire [62:0] _GEN_514 = {RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[
    31],RW0_wmask[30],_GEN_498};
  wire [63:0] _GEN_515 = {RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[31],RW0_wmask[
    31],RW0_wmask[31],RW0_wmask[30],_GEN_498};
  ip224uhdlp1p11rf_512x64m4b2c1s1_t0r0p0d0a1m1h mem_0_0 (
    .adr(mem_0_0_adr),
    .clk(mem_0_0_clk),
    .din(mem_0_0_din),
    .q(mem_0_0_q),
    .ren(mem_0_0_ren),
    .wen(mem_0_0_wen),
    .wbeb(mem_0_0_wbeb),
    .mcen(mem_0_0_mcen),
    .mc(mem_0_0_mc),
    .wa(mem_0_0_wa),
    .wpulse(mem_0_0_wpulse),
    .wpulseen(mem_0_0_wpulseen),
    .fwen(mem_0_0_fwen),
    .clkbyp(mem_0_0_clkbyp)
  );
  ip224uhdlp1p11rf_512x64m4b2c1s1_t0r0p0d0a1m1h mem_0_1 (
    .adr(mem_0_1_adr),
    .clk(mem_0_1_clk),
    .din(mem_0_1_din),
    .q(mem_0_1_q),
    .ren(mem_0_1_ren),
    .wen(mem_0_1_wen),
    .wbeb(mem_0_1_wbeb),
    .mcen(mem_0_1_mcen),
    .mc(mem_0_1_mc),
    .wa(mem_0_1_wa),
    .wpulse(mem_0_1_wpulse),
    .wpulseen(mem_0_1_wpulseen),
    .fwen(mem_0_1_fwen),
    .clkbyp(mem_0_1_clkbyp)
  );
  ip224uhdlp1p11rf_512x64m4b2c1s1_t0r0p0d0a1m1h mem_0_2 (
    .adr(mem_0_2_adr),
    .clk(mem_0_2_clk),
    .din(mem_0_2_din),
    .q(mem_0_2_q),
    .ren(mem_0_2_ren),
    .wen(mem_0_2_wen),
    .wbeb(mem_0_2_wbeb),
    .mcen(mem_0_2_mcen),
    .mc(mem_0_2_mc),
    .wa(mem_0_2_wa),
    .wpulse(mem_0_2_wpulse),
    .wpulseen(mem_0_2_wpulseen),
    .fwen(mem_0_2_fwen),
    .clkbyp(mem_0_2_clkbyp)
  );
  ip224uhdlp1p11rf_512x64m4b2c1s1_t0r0p0d0a1m1h mem_0_3 (
    .adr(mem_0_3_adr),
    .clk(mem_0_3_clk),
    .din(mem_0_3_din),
    .q(mem_0_3_q),
    .ren(mem_0_3_ren),
    .wen(mem_0_3_wen),
    .wbeb(mem_0_3_wbeb),
    .mcen(mem_0_3_mcen),
    .mc(mem_0_3_mc),
    .wa(mem_0_3_wa),
    .wpulse(mem_0_3_wpulse),
    .wpulseen(mem_0_3_wpulseen),
    .fwen(mem_0_3_fwen),
    .clkbyp(mem_0_3_clkbyp)
  );
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1};
  assign mem_0_0_adr = RW0_addr;
  assign mem_0_0_clk = RW0_clk;
  assign mem_0_0_din = RW0_wdata[63:0];
  assign mem_0_0_ren = ~RW0_wmode & RW0_en;
  assign mem_0_0_wen = RW0_wmode & RW0_en;
  assign mem_0_0_wbeb = ~_GEN_131;
  assign mem_0_0_mcen = 1'h0;
  assign mem_0_0_mc = 3'h0;
  assign mem_0_0_wa = 2'h0;
  assign mem_0_0_wpulse = 2'h0;
  assign mem_0_0_wpulseen = 1'h1;
  assign mem_0_0_fwen = 1'h0;
  assign mem_0_0_clkbyp = 1'h0;
  assign mem_0_1_adr = RW0_addr;
  assign mem_0_1_clk = RW0_clk;
  assign mem_0_1_din = RW0_wdata[127:64];
  assign mem_0_1_ren = ~RW0_wmode & RW0_en;
  assign mem_0_1_wen = RW0_wmode & RW0_en;
  assign mem_0_1_wbeb = ~_GEN_259;
  assign mem_0_1_mcen = 1'h0;
  assign mem_0_1_mc = 3'h0;
  assign mem_0_1_wa = 2'h0;
  assign mem_0_1_wpulse = 2'h0;
  assign mem_0_1_wpulseen = 1'h1;
  assign mem_0_1_fwen = 1'h0;
  assign mem_0_1_clkbyp = 1'h0;
  assign mem_0_2_adr = RW0_addr;
  assign mem_0_2_clk = RW0_clk;
  assign mem_0_2_din = RW0_wdata[191:128];
  assign mem_0_2_ren = ~RW0_wmode & RW0_en;
  assign mem_0_2_wen = RW0_wmode & RW0_en;
  assign mem_0_2_wbeb = ~_GEN_387;
  assign mem_0_2_mcen = 1'h0;
  assign mem_0_2_mc = 3'h0;
  assign mem_0_2_wa = 2'h0;
  assign mem_0_2_wpulse = 2'h0;
  assign mem_0_2_wpulseen = 1'h1;
  assign mem_0_2_fwen = 1'h0;
  assign mem_0_2_clkbyp = 1'h0;
  assign mem_0_3_adr = RW0_addr;
  assign mem_0_3_clk = RW0_clk;
  assign mem_0_3_din = RW0_wdata[255:192];
  assign mem_0_3_ren = ~RW0_wmode & RW0_en;
  assign mem_0_3_wen = RW0_wmode & RW0_en;
  assign mem_0_3_wbeb = ~_GEN_515;
  assign mem_0_3_mcen = 1'h0;
  assign mem_0_3_mc = 3'h0;
  assign mem_0_3_wa = 2'h0;
  assign mem_0_3_wpulse = 2'h0;
  assign mem_0_3_wpulseen = 1'h1;
  assign mem_0_3_fwen = 1'h0;
  assign mem_0_3_clkbyp = 1'h0;
endmodule
module tag_array_ext(
  input  [5:0]  RW0_addr,
  input         RW0_clk,
  input  [99:0] RW0_wdata,
  output [99:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input  [3:0]  RW0_wmask
);
  wire [8:0] mem_0_0_adr;
  wire  mem_0_0_clk;
  wire [49:0] mem_0_0_din;
  wire [49:0] mem_0_0_q;
  wire  mem_0_0_ren;
  wire  mem_0_0_wen;
  wire [49:0] mem_0_0_wbeb;
  wire  mem_0_0_mcen;
  wire [2:0] mem_0_0_mc;
  wire [1:0] mem_0_0_wa;
  wire [1:0] mem_0_0_wpulse;
  wire  mem_0_0_wpulseen;
  wire  mem_0_0_fwen;
  wire  mem_0_0_clkbyp;
  wire [8:0] mem_0_1_adr;
  wire  mem_0_1_clk;
  wire [49:0] mem_0_1_din;
  wire [49:0] mem_0_1_q;
  wire  mem_0_1_ren;
  wire  mem_0_1_wen;
  wire [49:0] mem_0_1_wbeb;
  wire  mem_0_1_mcen;
  wire [2:0] mem_0_1_mc;
  wire [1:0] mem_0_1_wa;
  wire [1:0] mem_0_1_wpulse;
  wire  mem_0_1_wpulseen;
  wire  mem_0_1_fwen;
  wire  mem_0_1_clkbyp;
  wire [49:0] RW0_rdata_0_0 = mem_0_0_q;
  wire [49:0] RW0_rdata_0_1 = mem_0_1_q;
  wire [99:0] RW0_rdata_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = RW0_wmask[0];
  wire  _GEN_2 = RW0_wmask[0];
  wire  _GEN_3 = RW0_wmask[0];
  wire [1:0] _GEN_4 = {RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_5 = RW0_wmask[0];
  wire [2:0] _GEN_6 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_7 = RW0_wmask[0];
  wire [3:0] _GEN_8 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_9 = RW0_wmask[0];
  wire [4:0] _GEN_10 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_11 = RW0_wmask[0];
  wire [5:0] _GEN_12 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_13 = RW0_wmask[0];
  wire [6:0] _GEN_14 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_15 = RW0_wmask[0];
  wire [7:0] _GEN_16 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0]};
  wire  _GEN_17 = RW0_wmask[0];
  wire [8:0] _GEN_18 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_19 = RW0_wmask[0];
  wire [9:0] _GEN_20 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_21 = RW0_wmask[0];
  wire [10:0] _GEN_22 = {RW0_wmask[0],_GEN_20};
  wire  _GEN_23 = RW0_wmask[0];
  wire [11:0] _GEN_24 = {RW0_wmask[0],RW0_wmask[0],_GEN_20};
  wire  _GEN_25 = RW0_wmask[0];
  wire [12:0] _GEN_26 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_20};
  wire  _GEN_27 = RW0_wmask[0];
  wire [13:0] _GEN_28 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_20};
  wire  _GEN_29 = RW0_wmask[0];
  wire [14:0] _GEN_30 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_20};
  wire  _GEN_31 = RW0_wmask[0];
  wire [15:0] _GEN_32 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_20};
  wire  _GEN_33 = RW0_wmask[0];
  wire [16:0] _GEN_34 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    _GEN_20};
  wire  _GEN_35 = RW0_wmask[0];
  wire [17:0] _GEN_36 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],_GEN_20};
  wire  _GEN_37 = RW0_wmask[0];
  wire [18:0] _GEN_38 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0],_GEN_20};
  wire  _GEN_39 = RW0_wmask[0];
  wire [19:0] _GEN_40 = {RW0_wmask[0],_GEN_38};
  wire  _GEN_41 = RW0_wmask[0];
  wire [20:0] _GEN_42 = {RW0_wmask[0],RW0_wmask[0],_GEN_38};
  wire  _GEN_43 = RW0_wmask[0];
  wire [21:0] _GEN_44 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_38};
  wire  _GEN_45 = RW0_wmask[0];
  wire [22:0] _GEN_46 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_38};
  wire  _GEN_47 = RW0_wmask[0];
  wire [23:0] _GEN_48 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_38};
  wire  _GEN_49 = RW0_wmask[1];
  wire [24:0] _GEN_50 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_38};
  wire  _GEN_51 = RW0_wmask[1];
  wire [25:0] _GEN_52 = {RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    _GEN_38};
  wire  _GEN_53 = RW0_wmask[1];
  wire [26:0] _GEN_54 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],_GEN_38};
  wire  _GEN_55 = RW0_wmask[1];
  wire [27:0] _GEN_56 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0],_GEN_38};
  wire  _GEN_57 = RW0_wmask[1];
  wire [28:0] _GEN_58 = {RW0_wmask[1],_GEN_56};
  wire  _GEN_59 = RW0_wmask[1];
  wire [29:0] _GEN_60 = {RW0_wmask[1],RW0_wmask[1],_GEN_56};
  wire  _GEN_61 = RW0_wmask[1];
  wire [30:0] _GEN_62 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_56};
  wire  _GEN_63 = RW0_wmask[1];
  wire [31:0] _GEN_64 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_56};
  wire  _GEN_65 = RW0_wmask[1];
  wire [32:0] _GEN_66 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_56};
  wire  _GEN_67 = RW0_wmask[1];
  wire [33:0] _GEN_68 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_56};
  wire  _GEN_69 = RW0_wmask[1];
  wire [34:0] _GEN_70 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    _GEN_56};
  wire  _GEN_71 = RW0_wmask[1];
  wire [35:0] _GEN_72 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],_GEN_56};
  wire  _GEN_73 = RW0_wmask[1];
  wire [36:0] _GEN_74 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],RW0_wmask[1],_GEN_56};
  wire  _GEN_75 = RW0_wmask[1];
  wire [37:0] _GEN_76 = {RW0_wmask[1],_GEN_74};
  wire  _GEN_77 = RW0_wmask[1];
  wire [38:0] _GEN_78 = {RW0_wmask[1],RW0_wmask[1],_GEN_74};
  wire  _GEN_79 = RW0_wmask[1];
  wire [39:0] _GEN_80 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_74};
  wire  _GEN_81 = RW0_wmask[1];
  wire [40:0] _GEN_82 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_74};
  wire  _GEN_83 = RW0_wmask[1];
  wire [41:0] _GEN_84 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_74};
  wire  _GEN_85 = RW0_wmask[1];
  wire [42:0] _GEN_86 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_74};
  wire  _GEN_87 = RW0_wmask[1];
  wire [43:0] _GEN_88 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    _GEN_74};
  wire  _GEN_89 = RW0_wmask[1];
  wire [44:0] _GEN_90 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],_GEN_74};
  wire  _GEN_91 = RW0_wmask[1];
  wire [45:0] _GEN_92 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],RW0_wmask[1],_GEN_74};
  wire  _GEN_93 = RW0_wmask[1];
  wire [46:0] _GEN_94 = {RW0_wmask[1],_GEN_92};
  wire  _GEN_95 = RW0_wmask[1];
  wire [47:0] _GEN_96 = {RW0_wmask[1],RW0_wmask[1],_GEN_92};
  wire  _GEN_97 = RW0_wmask[1];
  wire [48:0] _GEN_98 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_92};
  wire [49:0] _GEN_99 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_92};
  wire  _GEN_100 = ~RW0_wmode;
  wire  _GEN_101 = RW0_wmask[2];
  wire  _GEN_102 = RW0_wmask[2];
  wire  _GEN_103 = RW0_wmask[2];
  wire [1:0] _GEN_104 = {RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_105 = RW0_wmask[2];
  wire [2:0] _GEN_106 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_107 = RW0_wmask[2];
  wire [3:0] _GEN_108 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_109 = RW0_wmask[2];
  wire [4:0] _GEN_110 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_111 = RW0_wmask[2];
  wire [5:0] _GEN_112 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_113 = RW0_wmask[2];
  wire [6:0] _GEN_114 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_115 = RW0_wmask[2];
  wire [7:0] _GEN_116 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2]};
  wire  _GEN_117 = RW0_wmask[2];
  wire [8:0] _GEN_118 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_119 = RW0_wmask[2];
  wire [9:0] _GEN_120 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_121 = RW0_wmask[2];
  wire [10:0] _GEN_122 = {RW0_wmask[2],_GEN_120};
  wire  _GEN_123 = RW0_wmask[2];
  wire [11:0] _GEN_124 = {RW0_wmask[2],RW0_wmask[2],_GEN_120};
  wire  _GEN_125 = RW0_wmask[2];
  wire [12:0] _GEN_126 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_120};
  wire  _GEN_127 = RW0_wmask[2];
  wire [13:0] _GEN_128 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_120};
  wire  _GEN_129 = RW0_wmask[2];
  wire [14:0] _GEN_130 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_120};
  wire  _GEN_131 = RW0_wmask[2];
  wire [15:0] _GEN_132 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_120};
  wire  _GEN_133 = RW0_wmask[2];
  wire [16:0] _GEN_134 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    _GEN_120};
  wire  _GEN_135 = RW0_wmask[2];
  wire [17:0] _GEN_136 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],_GEN_120};
  wire  _GEN_137 = RW0_wmask[2];
  wire [18:0] _GEN_138 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],RW0_wmask[2],_GEN_120};
  wire  _GEN_139 = RW0_wmask[2];
  wire [19:0] _GEN_140 = {RW0_wmask[2],_GEN_138};
  wire  _GEN_141 = RW0_wmask[2];
  wire [20:0] _GEN_142 = {RW0_wmask[2],RW0_wmask[2],_GEN_138};
  wire  _GEN_143 = RW0_wmask[2];
  wire [21:0] _GEN_144 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_138};
  wire  _GEN_145 = RW0_wmask[2];
  wire [22:0] _GEN_146 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_138};
  wire  _GEN_147 = RW0_wmask[2];
  wire [23:0] _GEN_148 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_138};
  wire  _GEN_149 = RW0_wmask[3];
  wire [24:0] _GEN_150 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_138};
  wire  _GEN_151 = RW0_wmask[3];
  wire [25:0] _GEN_152 = {RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    _GEN_138};
  wire  _GEN_153 = RW0_wmask[3];
  wire [26:0] _GEN_154 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],_GEN_138};
  wire  _GEN_155 = RW0_wmask[3];
  wire [27:0] _GEN_156 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],RW0_wmask[2],_GEN_138};
  wire  _GEN_157 = RW0_wmask[3];
  wire [28:0] _GEN_158 = {RW0_wmask[3],_GEN_156};
  wire  _GEN_159 = RW0_wmask[3];
  wire [29:0] _GEN_160 = {RW0_wmask[3],RW0_wmask[3],_GEN_156};
  wire  _GEN_161 = RW0_wmask[3];
  wire [30:0] _GEN_162 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_156};
  wire  _GEN_163 = RW0_wmask[3];
  wire [31:0] _GEN_164 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_156};
  wire  _GEN_165 = RW0_wmask[3];
  wire [32:0] _GEN_166 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_156};
  wire  _GEN_167 = RW0_wmask[3];
  wire [33:0] _GEN_168 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_156};
  wire  _GEN_169 = RW0_wmask[3];
  wire [34:0] _GEN_170 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    _GEN_156};
  wire  _GEN_171 = RW0_wmask[3];
  wire [35:0] _GEN_172 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],_GEN_156};
  wire  _GEN_173 = RW0_wmask[3];
  wire [36:0] _GEN_174 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],RW0_wmask[3],_GEN_156};
  wire  _GEN_175 = RW0_wmask[3];
  wire [37:0] _GEN_176 = {RW0_wmask[3],_GEN_174};
  wire  _GEN_177 = RW0_wmask[3];
  wire [38:0] _GEN_178 = {RW0_wmask[3],RW0_wmask[3],_GEN_174};
  wire  _GEN_179 = RW0_wmask[3];
  wire [39:0] _GEN_180 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_174};
  wire  _GEN_181 = RW0_wmask[3];
  wire [40:0] _GEN_182 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_174};
  wire  _GEN_183 = RW0_wmask[3];
  wire [41:0] _GEN_184 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_174};
  wire  _GEN_185 = RW0_wmask[3];
  wire [42:0] _GEN_186 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_174};
  wire  _GEN_187 = RW0_wmask[3];
  wire [43:0] _GEN_188 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    _GEN_174};
  wire  _GEN_189 = RW0_wmask[3];
  wire [44:0] _GEN_190 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],_GEN_174};
  wire  _GEN_191 = RW0_wmask[3];
  wire [45:0] _GEN_192 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],RW0_wmask[3],_GEN_174};
  wire  _GEN_193 = RW0_wmask[3];
  wire [46:0] _GEN_194 = {RW0_wmask[3],_GEN_192};
  wire  _GEN_195 = RW0_wmask[3];
  wire [47:0] _GEN_196 = {RW0_wmask[3],RW0_wmask[3],_GEN_192};
  wire  _GEN_197 = RW0_wmask[3];
  wire [48:0] _GEN_198 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_192};
  wire [49:0] _GEN_199 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_192};
  ip224uhdlp1p11rf_512x50m4b2c1s1_t0r0p0d0a1m1h mem_0_0 (
    .adr(mem_0_0_adr),
    .clk(mem_0_0_clk),
    .din(mem_0_0_din),
    .q(mem_0_0_q),
    .ren(mem_0_0_ren),
    .wen(mem_0_0_wen),
    .wbeb(mem_0_0_wbeb),
    .mcen(mem_0_0_mcen),
    .mc(mem_0_0_mc),
    .wa(mem_0_0_wa),
    .wpulse(mem_0_0_wpulse),
    .wpulseen(mem_0_0_wpulseen),
    .fwen(mem_0_0_fwen),
    .clkbyp(mem_0_0_clkbyp)
  );
  ip224uhdlp1p11rf_512x50m4b2c1s1_t0r0p0d0a1m1h mem_0_1 (
    .adr(mem_0_1_adr),
    .clk(mem_0_1_clk),
    .din(mem_0_1_din),
    .q(mem_0_1_q),
    .ren(mem_0_1_ren),
    .wen(mem_0_1_wen),
    .wbeb(mem_0_1_wbeb),
    .mcen(mem_0_1_mcen),
    .mc(mem_0_1_mc),
    .wa(mem_0_1_wa),
    .wpulse(mem_0_1_wpulse),
    .wpulseen(mem_0_1_wpulseen),
    .fwen(mem_0_1_fwen),
    .clkbyp(mem_0_1_clkbyp)
  );
  assign RW0_rdata = {RW0_rdata_0_1,RW0_rdata_0_0};
  assign mem_0_0_adr = {{3'd0}, RW0_addr};
  assign mem_0_0_clk = RW0_clk;
  assign mem_0_0_din = RW0_wdata[49:0];
  assign mem_0_0_ren = ~RW0_wmode & RW0_en;
  assign mem_0_0_wen = RW0_wmode & RW0_en;
  assign mem_0_0_wbeb = ~_GEN_99;
  assign mem_0_0_mcen = 1'h0;
  assign mem_0_0_mc = 3'h0;
  assign mem_0_0_wa = 2'h0;
  assign mem_0_0_wpulse = 2'h0;
  assign mem_0_0_wpulseen = 1'h1;
  assign mem_0_0_fwen = 1'h0;
  assign mem_0_0_clkbyp = 1'h0;
  assign mem_0_1_adr = {{3'd0}, RW0_addr};
  assign mem_0_1_clk = RW0_clk;
  assign mem_0_1_din = RW0_wdata[99:50];
  assign mem_0_1_ren = ~RW0_wmode & RW0_en;
  assign mem_0_1_wen = RW0_wmode & RW0_en;
  assign mem_0_1_wbeb = ~_GEN_199;
  assign mem_0_1_mcen = 1'h0;
  assign mem_0_1_mc = 3'h0;
  assign mem_0_1_wa = 2'h0;
  assign mem_0_1_wpulse = 2'h0;
  assign mem_0_1_wpulseen = 1'h1;
  assign mem_0_1_fwen = 1'h0;
  assign mem_0_1_clkbyp = 1'h0;
endmodule
module tag_array_0_ext(
  input  [5:0]  RW0_addr,
  input         RW0_clk,
  input  [23:0] RW0_wdata,
  output [23:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode
);
  wire [8:0] mem_0_0_adr;
  wire  mem_0_0_clk;
  wire [23:0] mem_0_0_din;
  wire [23:0] mem_0_0_q;
  wire  mem_0_0_ren;
  wire  mem_0_0_wen;
  wire  mem_0_0_mcen;
  wire [2:0] mem_0_0_mc;
  wire [1:0] mem_0_0_wa;
  wire [1:0] mem_0_0_wpulse;
  wire  mem_0_0_wpulseen;
  wire  mem_0_0_fwen;
  wire  mem_0_0_clkbyp;
  wire [23:0] RW0_rdata_0_0 = mem_0_0_q;
  wire [23:0] RW0_rdata_0 = RW0_rdata_0_0;
  wire  _GEN_0 = ~RW0_wmode;
  ip224uhdlp1p11rf_512x24m4b2c1s0_t0r0p0d0a1m1h mem_0_0 (
    .adr(mem_0_0_adr),
    .clk(mem_0_0_clk),
    .din(mem_0_0_din),
    .q(mem_0_0_q),
    .ren(mem_0_0_ren),
    .wen(mem_0_0_wen),
    .mcen(mem_0_0_mcen),
    .mc(mem_0_0_mc),
    .wa(mem_0_0_wa),
    .wpulse(mem_0_0_wpulse),
    .wpulseen(mem_0_0_wpulseen),
    .fwen(mem_0_0_fwen),
    .clkbyp(mem_0_0_clkbyp)
  );
  assign RW0_rdata = mem_0_0_q;
  assign mem_0_0_adr = {{3'd0}, RW0_addr};
  assign mem_0_0_clk = RW0_clk;
  assign mem_0_0_din = RW0_wdata;
  assign mem_0_0_ren = ~RW0_wmode & RW0_en;
  assign mem_0_0_wen = RW0_wmode & RW0_en;
  assign mem_0_0_mcen = 1'h0;
  assign mem_0_0_mc = 3'h0;
  assign mem_0_0_wa = 2'h0;
  assign mem_0_0_wpulse = 2'h0;
  assign mem_0_0_wpulseen = 1'h1;
  assign mem_0_0_fwen = 1'h0;
  assign mem_0_0_clkbyp = 1'h0;
endmodule
module data_arrays_0_0_ext(
  input  [8:0]  RW0_addr,
  input         RW0_clk,
  input  [31:0] RW0_wdata,
  output [31:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode
);
  wire [8:0] mem_0_0_adr;
  wire  mem_0_0_clk;
  wire [31:0] mem_0_0_din;
  wire [31:0] mem_0_0_q;
  wire  mem_0_0_ren;
  wire  mem_0_0_wen;
  wire  mem_0_0_mcen;
  wire [2:0] mem_0_0_mc;
  wire [1:0] mem_0_0_wa;
  wire [1:0] mem_0_0_wpulse;
  wire  mem_0_0_wpulseen;
  wire  mem_0_0_fwen;
  wire  mem_0_0_clkbyp;
  wire [31:0] RW0_rdata_0_0 = mem_0_0_q;
  wire [31:0] RW0_rdata_0 = RW0_rdata_0_0;
  wire  _GEN_0 = ~RW0_wmode;
  ip224uhdlp1p11rf_512x32m4b2c1s0_t0r0p0d0a1m1h mem_0_0 (
    .adr(mem_0_0_adr),
    .clk(mem_0_0_clk),
    .din(mem_0_0_din),
    .q(mem_0_0_q),
    .ren(mem_0_0_ren),
    .wen(mem_0_0_wen),
    .mcen(mem_0_0_mcen),
    .mc(mem_0_0_mc),
    .wa(mem_0_0_wa),
    .wpulse(mem_0_0_wpulse),
    .wpulseen(mem_0_0_wpulseen),
    .fwen(mem_0_0_fwen),
    .clkbyp(mem_0_0_clkbyp)
  );
  assign RW0_rdata = mem_0_0_q;
  assign mem_0_0_adr = RW0_addr;
  assign mem_0_0_clk = RW0_clk;
  assign mem_0_0_din = RW0_wdata;
  assign mem_0_0_ren = ~RW0_wmode & RW0_en;
  assign mem_0_0_wen = RW0_wmode & RW0_en;
  assign mem_0_0_mcen = 1'h0;
  assign mem_0_0_mc = 3'h0;
  assign mem_0_0_wa = 2'h0;
  assign mem_0_0_wpulse = 2'h0;
  assign mem_0_0_wpulseen = 1'h1;
  assign mem_0_0_fwen = 1'h0;
  assign mem_0_0_clkbyp = 1'h0;
endmodule
module tag_array_1_ext(
  input  [5:0]  R0_addr,
  input         R0_clk,
  output [99:0] R0_data,
  input         R0_en,
  input  [5:0]  W0_addr,
  input         W0_clk,
  input  [99:0] W0_data,
  input         W0_en,
  input  [3:0]  W0_mask
);
  wire [5:0] mem_0_0_iarp0;
  wire  mem_0_0_ickrp0;
  wire [99:0] mem_0_0_odoutp0;
  wire  mem_0_0_irenp0;
  wire [5:0] mem_0_0_iawp0;
  wire  mem_0_0_ickwp0;
  wire [99:0] mem_0_0_idinp0;
  wire  mem_0_0_iwenp0;
  wire [99:0] mem_0_0_ibwep0;
  wire  mem_0_0_ifuse;
  wire  mem_0_0_iclkbyp;
  wire  mem_0_0_imce;
  wire [1:0] mem_0_0_irmce;
  wire [3:0] mem_0_0_iwmce;
  wire [99:0] R0_data_0_0 = mem_0_0_odoutp0;
  wire [99:0] R0_data_0 = R0_data_0_0;
  wire  _GEN_0 = W0_mask[0];
  wire  _GEN_1 = W0_mask[0];
  wire  _GEN_2 = W0_mask[0];
  wire [1:0] _GEN_3 = {W0_mask[0],W0_mask[0]};
  wire  _GEN_4 = W0_mask[0];
  wire [2:0] _GEN_5 = {W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_6 = W0_mask[0];
  wire [3:0] _GEN_7 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_8 = W0_mask[0];
  wire [4:0] _GEN_9 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_10 = W0_mask[0];
  wire [5:0] _GEN_11 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_12 = W0_mask[0];
  wire [6:0] _GEN_13 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_14 = W0_mask[0];
  wire [7:0] _GEN_15 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_16 = W0_mask[0];
  wire [8:0] _GEN_17 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[
    0]};
  wire  _GEN_18 = W0_mask[0];
  wire [9:0] _GEN_19 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[
    0],W0_mask[0]};
  wire  _GEN_20 = W0_mask[0];
  wire [10:0] _GEN_21 = {W0_mask[0],_GEN_19};
  wire  _GEN_22 = W0_mask[0];
  wire [11:0] _GEN_23 = {W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_24 = W0_mask[0];
  wire [12:0] _GEN_25 = {W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_26 = W0_mask[0];
  wire [13:0] _GEN_27 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_28 = W0_mask[0];
  wire [14:0] _GEN_29 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_30 = W0_mask[0];
  wire [15:0] _GEN_31 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_32 = W0_mask[0];
  wire [16:0] _GEN_33 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_34 = W0_mask[0];
  wire [17:0] _GEN_35 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19
    };
  wire  _GEN_36 = W0_mask[0];
  wire [18:0] _GEN_37 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask
    [0],_GEN_19};
  wire  _GEN_38 = W0_mask[0];
  wire [19:0] _GEN_39 = {W0_mask[0],_GEN_37};
  wire  _GEN_40 = W0_mask[0];
  wire [20:0] _GEN_41 = {W0_mask[0],W0_mask[0],_GEN_37};
  wire  _GEN_42 = W0_mask[0];
  wire [21:0] _GEN_43 = {W0_mask[0],W0_mask[0],W0_mask[0],_GEN_37};
  wire  _GEN_44 = W0_mask[0];
  wire [22:0] _GEN_45 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_37};
  wire  _GEN_46 = W0_mask[0];
  wire [23:0] _GEN_47 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_37};
  wire  _GEN_48 = W0_mask[1];
  wire [24:0] _GEN_49 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_37};
  wire  _GEN_50 = W0_mask[1];
  wire [25:0] _GEN_51 = {W0_mask[1],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_37};
  wire  _GEN_52 = W0_mask[1];
  wire [26:0] _GEN_53 = {W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_37
    };
  wire  _GEN_54 = W0_mask[1];
  wire [27:0] _GEN_55 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask
    [0],_GEN_37};
  wire  _GEN_56 = W0_mask[1];
  wire [28:0] _GEN_57 = {W0_mask[1],_GEN_55};
  wire  _GEN_58 = W0_mask[1];
  wire [29:0] _GEN_59 = {W0_mask[1],W0_mask[1],_GEN_55};
  wire  _GEN_60 = W0_mask[1];
  wire [30:0] _GEN_61 = {W0_mask[1],W0_mask[1],W0_mask[1],_GEN_55};
  wire  _GEN_62 = W0_mask[1];
  wire [31:0] _GEN_63 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_55};
  wire  _GEN_64 = W0_mask[1];
  wire [32:0] _GEN_65 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_55};
  wire  _GEN_66 = W0_mask[1];
  wire [33:0] _GEN_67 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_55};
  wire  _GEN_68 = W0_mask[1];
  wire [34:0] _GEN_69 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_55};
  wire  _GEN_70 = W0_mask[1];
  wire [35:0] _GEN_71 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_55
    };
  wire  _GEN_72 = W0_mask[1];
  wire [36:0] _GEN_73 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask
    [1],_GEN_55};
  wire  _GEN_74 = W0_mask[1];
  wire [37:0] _GEN_75 = {W0_mask[1],_GEN_73};
  wire  _GEN_76 = W0_mask[1];
  wire [38:0] _GEN_77 = {W0_mask[1],W0_mask[1],_GEN_73};
  wire  _GEN_78 = W0_mask[1];
  wire [39:0] _GEN_79 = {W0_mask[1],W0_mask[1],W0_mask[1],_GEN_73};
  wire  _GEN_80 = W0_mask[1];
  wire [40:0] _GEN_81 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_73};
  wire  _GEN_82 = W0_mask[1];
  wire [41:0] _GEN_83 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_73};
  wire  _GEN_84 = W0_mask[1];
  wire [42:0] _GEN_85 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_73};
  wire  _GEN_86 = W0_mask[1];
  wire [43:0] _GEN_87 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_73};
  wire  _GEN_88 = W0_mask[1];
  wire [44:0] _GEN_89 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_73
    };
  wire  _GEN_90 = W0_mask[1];
  wire [45:0] _GEN_91 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask
    [1],_GEN_73};
  wire  _GEN_92 = W0_mask[1];
  wire [46:0] _GEN_93 = {W0_mask[1],_GEN_91};
  wire  _GEN_94 = W0_mask[1];
  wire [47:0] _GEN_95 = {W0_mask[1],W0_mask[1],_GEN_91};
  wire  _GEN_96 = W0_mask[1];
  wire [48:0] _GEN_97 = {W0_mask[1],W0_mask[1],W0_mask[1],_GEN_91};
  wire  _GEN_98 = W0_mask[2];
  wire [49:0] _GEN_99 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_91};
  wire  _GEN_100 = W0_mask[2];
  wire [50:0] _GEN_101 = {W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_91};
  wire  _GEN_102 = W0_mask[2];
  wire [51:0] _GEN_103 = {W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_91};
  wire  _GEN_104 = W0_mask[2];
  wire [52:0] _GEN_105 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_91};
  wire  _GEN_106 = W0_mask[2];
  wire [53:0] _GEN_107 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],
    _GEN_91};
  wire  _GEN_108 = W0_mask[2];
  wire [54:0] _GEN_109 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],
    W0_mask[1],_GEN_91};
  wire  _GEN_110 = W0_mask[2];
  wire [55:0] _GEN_111 = {W0_mask[2],_GEN_109};
  wire  _GEN_112 = W0_mask[2];
  wire [56:0] _GEN_113 = {W0_mask[2],W0_mask[2],_GEN_109};
  wire  _GEN_114 = W0_mask[2];
  wire [57:0] _GEN_115 = {W0_mask[2],W0_mask[2],W0_mask[2],_GEN_109};
  wire  _GEN_116 = W0_mask[2];
  wire [58:0] _GEN_117 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_109};
  wire  _GEN_118 = W0_mask[2];
  wire [59:0] _GEN_119 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_109};
  wire  _GEN_120 = W0_mask[2];
  wire [60:0] _GEN_121 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_109};
  wire  _GEN_122 = W0_mask[2];
  wire [61:0] _GEN_123 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_109};
  wire  _GEN_124 = W0_mask[2];
  wire [62:0] _GEN_125 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],
    _GEN_109};
  wire  _GEN_126 = W0_mask[2];
  wire [63:0] _GEN_127 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],
    W0_mask[2],_GEN_109};
  wire  _GEN_128 = W0_mask[2];
  wire [64:0] _GEN_129 = {W0_mask[2],_GEN_127};
  wire  _GEN_130 = W0_mask[2];
  wire [65:0] _GEN_131 = {W0_mask[2],W0_mask[2],_GEN_127};
  wire  _GEN_132 = W0_mask[2];
  wire [66:0] _GEN_133 = {W0_mask[2],W0_mask[2],W0_mask[2],_GEN_127};
  wire  _GEN_134 = W0_mask[2];
  wire [67:0] _GEN_135 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_127};
  wire  _GEN_136 = W0_mask[2];
  wire [68:0] _GEN_137 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_127};
  wire  _GEN_138 = W0_mask[2];
  wire [69:0] _GEN_139 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_127};
  wire  _GEN_140 = W0_mask[2];
  wire [70:0] _GEN_141 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_127};
  wire  _GEN_142 = W0_mask[2];
  wire [71:0] _GEN_143 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],
    _GEN_127};
  wire  _GEN_144 = W0_mask[2];
  wire [72:0] _GEN_145 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],
    W0_mask[2],_GEN_127};
  wire  _GEN_146 = W0_mask[2];
  wire [73:0] _GEN_147 = {W0_mask[2],_GEN_145};
  wire  _GEN_148 = W0_mask[3];
  wire [74:0] _GEN_149 = {W0_mask[2],W0_mask[2],_GEN_145};
  wire  _GEN_150 = W0_mask[3];
  wire [75:0] _GEN_151 = {W0_mask[3],W0_mask[2],W0_mask[2],_GEN_145};
  wire  _GEN_152 = W0_mask[3];
  wire [76:0] _GEN_153 = {W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],_GEN_145};
  wire  _GEN_154 = W0_mask[3];
  wire [77:0] _GEN_155 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],_GEN_145};
  wire  _GEN_156 = W0_mask[3];
  wire [78:0] _GEN_157 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],_GEN_145};
  wire  _GEN_158 = W0_mask[3];
  wire [79:0] _GEN_159 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],_GEN_145};
  wire  _GEN_160 = W0_mask[3];
  wire [80:0] _GEN_161 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],
    _GEN_145};
  wire  _GEN_162 = W0_mask[3];
  wire [81:0] _GEN_163 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],
    W0_mask[2],_GEN_145};
  wire  _GEN_164 = W0_mask[3];
  wire [82:0] _GEN_165 = {W0_mask[3],_GEN_163};
  wire  _GEN_166 = W0_mask[3];
  wire [83:0] _GEN_167 = {W0_mask[3],W0_mask[3],_GEN_163};
  wire  _GEN_168 = W0_mask[3];
  wire [84:0] _GEN_169 = {W0_mask[3],W0_mask[3],W0_mask[3],_GEN_163};
  wire  _GEN_170 = W0_mask[3];
  wire [85:0] _GEN_171 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_163};
  wire  _GEN_172 = W0_mask[3];
  wire [86:0] _GEN_173 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_163};
  wire  _GEN_174 = W0_mask[3];
  wire [87:0] _GEN_175 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_163};
  wire  _GEN_176 = W0_mask[3];
  wire [88:0] _GEN_177 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_163};
  wire  _GEN_178 = W0_mask[3];
  wire [89:0] _GEN_179 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],
    _GEN_163};
  wire  _GEN_180 = W0_mask[3];
  wire [90:0] _GEN_181 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],
    W0_mask[3],_GEN_163};
  wire  _GEN_182 = W0_mask[3];
  wire [91:0] _GEN_183 = {W0_mask[3],_GEN_181};
  wire  _GEN_184 = W0_mask[3];
  wire [92:0] _GEN_185 = {W0_mask[3],W0_mask[3],_GEN_181};
  wire  _GEN_186 = W0_mask[3];
  wire [93:0] _GEN_187 = {W0_mask[3],W0_mask[3],W0_mask[3],_GEN_181};
  wire  _GEN_188 = W0_mask[3];
  wire [94:0] _GEN_189 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_181};
  wire  _GEN_190 = W0_mask[3];
  wire [95:0] _GEN_191 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_181};
  wire  _GEN_192 = W0_mask[3];
  wire [96:0] _GEN_193 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_181};
  wire  _GEN_194 = W0_mask[3];
  wire [97:0] _GEN_195 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_181};
  wire  _GEN_196 = W0_mask[3];
  wire [98:0] _GEN_197 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],
    _GEN_181};
  ip224rfsbhpm1r1w64x100be100m1 mem_0_0 (
    .iarp0(mem_0_0_iarp0),
    .ickrp0(mem_0_0_ickrp0),
    .odoutp0(mem_0_0_odoutp0),
    .irenp0(mem_0_0_irenp0),
    .iawp0(mem_0_0_iawp0),
    .ickwp0(mem_0_0_ickwp0),
    .idinp0(mem_0_0_idinp0),
    .iwenp0(mem_0_0_iwenp0),
    .ibwep0(mem_0_0_ibwep0),
    .ifuse(mem_0_0_ifuse),
    .iclkbyp(mem_0_0_iclkbyp),
    .imce(mem_0_0_imce),
    .irmce(mem_0_0_irmce),
    .iwmce(mem_0_0_iwmce)
  );
  assign R0_data = mem_0_0_odoutp0;
  assign mem_0_0_iarp0 = R0_addr;
  assign mem_0_0_ickrp0 = R0_clk;
  assign mem_0_0_irenp0 = R0_en;
  assign mem_0_0_iawp0 = W0_addr;
  assign mem_0_0_ickwp0 = W0_clk;
  assign mem_0_0_idinp0 = W0_data;
  assign mem_0_0_iwenp0 = W0_en;
  assign mem_0_0_ibwep0 = {W0_mask[3],_GEN_197};
  assign mem_0_0_ifuse = 1'h0;
  assign mem_0_0_iclkbyp = 1'h0;
  assign mem_0_0_imce = 1'h0;
  assign mem_0_0_irmce = 2'h0;
  assign mem_0_0_iwmce = 4'h0;
endmodule
module array_0_0_0_ext(
  input  [8:0]  R0_addr,
  input         R0_clk,
  output [63:0] R0_data,
  input         R0_en,
  input  [8:0]  W0_addr,
  input         W0_clk,
  input  [63:0] W0_data,
  input         W0_en
);
  wire [8:0] mem_0_0_iarp0;
  wire  mem_0_0_ickrp0;
  wire [63:0] mem_0_0_odoutp0;
  wire  mem_0_0_irenp0;
  wire [8:0] mem_0_0_iawp0;
  wire  mem_0_0_ickwp0;
  wire [63:0] mem_0_0_idinp0;
  wire  mem_0_0_iwenp0;
  wire  mem_0_0_ifuse;
  wire  mem_0_0_iclkbyp;
  wire  mem_0_0_imce;
  wire [1:0] mem_0_0_irmce;
  wire [3:0] mem_0_0_iwmce;
  wire [63:0] R0_data_0_0 = mem_0_0_odoutp0;
  wire [63:0] R0_data_0 = R0_data_0_0;
  ip224rfsbhpm1r1w512x64m1 mem_0_0 (
    .iarp0(mem_0_0_iarp0),
    .ickrp0(mem_0_0_ickrp0),
    .odoutp0(mem_0_0_odoutp0),
    .irenp0(mem_0_0_irenp0),
    .iawp0(mem_0_0_iawp0),
    .ickwp0(mem_0_0_ickwp0),
    .idinp0(mem_0_0_idinp0),
    .iwenp0(mem_0_0_iwenp0),
    .ifuse(mem_0_0_ifuse),
    .iclkbyp(mem_0_0_iclkbyp),
    .imce(mem_0_0_imce),
    .irmce(mem_0_0_irmce),
    .iwmce(mem_0_0_iwmce)
  );
  assign R0_data = mem_0_0_odoutp0;
  assign mem_0_0_iarp0 = R0_addr;
  assign mem_0_0_ickrp0 = R0_clk;
  assign mem_0_0_irenp0 = R0_en;
  assign mem_0_0_iawp0 = W0_addr;
  assign mem_0_0_ickwp0 = W0_clk;
  assign mem_0_0_idinp0 = W0_data;
  assign mem_0_0_iwenp0 = W0_en;
  assign mem_0_0_ifuse = 1'h0;
  assign mem_0_0_iclkbyp = 1'h0;
  assign mem_0_0_imce = 1'h0;
  assign mem_0_0_irmce = 2'h0;
  assign mem_0_0_iwmce = 4'h0;
endmodule
module tag_array_2_ext(
  input  [5:0]  RW0_addr,
  input         RW0_clk,
  input  [91:0] RW0_wdata,
  output [91:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input  [3:0]  RW0_wmask
);
  wire [8:0] mem_0_0_adr;
  wire  mem_0_0_clk;
  wire [45:0] mem_0_0_din;
  wire [45:0] mem_0_0_q;
  wire  mem_0_0_ren;
  wire  mem_0_0_wen;
  wire [45:0] mem_0_0_wbeb;
  wire  mem_0_0_mcen;
  wire [2:0] mem_0_0_mc;
  wire [1:0] mem_0_0_wa;
  wire [1:0] mem_0_0_wpulse;
  wire  mem_0_0_wpulseen;
  wire  mem_0_0_fwen;
  wire  mem_0_0_clkbyp;
  wire [8:0] mem_0_1_adr;
  wire  mem_0_1_clk;
  wire [45:0] mem_0_1_din;
  wire [45:0] mem_0_1_q;
  wire  mem_0_1_ren;
  wire  mem_0_1_wen;
  wire [45:0] mem_0_1_wbeb;
  wire  mem_0_1_mcen;
  wire [2:0] mem_0_1_mc;
  wire [1:0] mem_0_1_wa;
  wire [1:0] mem_0_1_wpulse;
  wire  mem_0_1_wpulseen;
  wire  mem_0_1_fwen;
  wire  mem_0_1_clkbyp;
  wire [45:0] RW0_rdata_0_0 = mem_0_0_q;
  wire [45:0] RW0_rdata_0_1 = mem_0_1_q;
  wire [91:0] RW0_rdata_0 = {RW0_rdata_0_1,RW0_rdata_0_0};
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = RW0_wmask[0];
  wire  _GEN_2 = RW0_wmask[0];
  wire  _GEN_3 = RW0_wmask[0];
  wire [1:0] _GEN_4 = {RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_5 = RW0_wmask[0];
  wire [2:0] _GEN_6 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_7 = RW0_wmask[0];
  wire [3:0] _GEN_8 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_9 = RW0_wmask[0];
  wire [4:0] _GEN_10 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_11 = RW0_wmask[0];
  wire [5:0] _GEN_12 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_13 = RW0_wmask[0];
  wire [6:0] _GEN_14 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_15 = RW0_wmask[0];
  wire [7:0] _GEN_16 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0]};
  wire  _GEN_17 = RW0_wmask[0];
  wire [8:0] _GEN_18 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_19 = RW0_wmask[0];
  wire [9:0] _GEN_20 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0],RW0_wmask[0]};
  wire  _GEN_21 = RW0_wmask[0];
  wire [10:0] _GEN_22 = {RW0_wmask[0],_GEN_20};
  wire  _GEN_23 = RW0_wmask[0];
  wire [11:0] _GEN_24 = {RW0_wmask[0],RW0_wmask[0],_GEN_20};
  wire  _GEN_25 = RW0_wmask[0];
  wire [12:0] _GEN_26 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_20};
  wire  _GEN_27 = RW0_wmask[0];
  wire [13:0] _GEN_28 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_20};
  wire  _GEN_29 = RW0_wmask[0];
  wire [14:0] _GEN_30 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_20};
  wire  _GEN_31 = RW0_wmask[0];
  wire [15:0] _GEN_32 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_20};
  wire  _GEN_33 = RW0_wmask[0];
  wire [16:0] _GEN_34 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    _GEN_20};
  wire  _GEN_35 = RW0_wmask[0];
  wire [17:0] _GEN_36 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],_GEN_20};
  wire  _GEN_37 = RW0_wmask[0];
  wire [18:0] _GEN_38 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0],_GEN_20};
  wire  _GEN_39 = RW0_wmask[0];
  wire [19:0] _GEN_40 = {RW0_wmask[0],_GEN_38};
  wire  _GEN_41 = RW0_wmask[0];
  wire [20:0] _GEN_42 = {RW0_wmask[0],RW0_wmask[0],_GEN_38};
  wire  _GEN_43 = RW0_wmask[0];
  wire [21:0] _GEN_44 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_38};
  wire  _GEN_45 = RW0_wmask[1];
  wire [22:0] _GEN_46 = {RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_38};
  wire  _GEN_47 = RW0_wmask[1];
  wire [23:0] _GEN_48 = {RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_38};
  wire  _GEN_49 = RW0_wmask[1];
  wire [24:0] _GEN_50 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],_GEN_38};
  wire  _GEN_51 = RW0_wmask[1];
  wire [25:0] _GEN_52 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    _GEN_38};
  wire  _GEN_53 = RW0_wmask[1];
  wire [26:0] _GEN_54 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],_GEN_38};
  wire  _GEN_55 = RW0_wmask[1];
  wire [27:0] _GEN_56 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[0],RW0_wmask[0],
    RW0_wmask[0],RW0_wmask[0],_GEN_38};
  wire  _GEN_57 = RW0_wmask[1];
  wire [28:0] _GEN_58 = {RW0_wmask[1],_GEN_56};
  wire  _GEN_59 = RW0_wmask[1];
  wire [29:0] _GEN_60 = {RW0_wmask[1],RW0_wmask[1],_GEN_56};
  wire  _GEN_61 = RW0_wmask[1];
  wire [30:0] _GEN_62 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_56};
  wire  _GEN_63 = RW0_wmask[1];
  wire [31:0] _GEN_64 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_56};
  wire  _GEN_65 = RW0_wmask[1];
  wire [32:0] _GEN_66 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_56};
  wire  _GEN_67 = RW0_wmask[1];
  wire [33:0] _GEN_68 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_56};
  wire  _GEN_69 = RW0_wmask[1];
  wire [34:0] _GEN_70 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    _GEN_56};
  wire  _GEN_71 = RW0_wmask[1];
  wire [35:0] _GEN_72 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],_GEN_56};
  wire  _GEN_73 = RW0_wmask[1];
  wire [36:0] _GEN_74 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],RW0_wmask[1],_GEN_56};
  wire  _GEN_75 = RW0_wmask[1];
  wire [37:0] _GEN_76 = {RW0_wmask[1],_GEN_74};
  wire  _GEN_77 = RW0_wmask[1];
  wire [38:0] _GEN_78 = {RW0_wmask[1],RW0_wmask[1],_GEN_74};
  wire  _GEN_79 = RW0_wmask[1];
  wire [39:0] _GEN_80 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_74};
  wire  _GEN_81 = RW0_wmask[1];
  wire [40:0] _GEN_82 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_74};
  wire  _GEN_83 = RW0_wmask[1];
  wire [41:0] _GEN_84 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_74};
  wire  _GEN_85 = RW0_wmask[1];
  wire [42:0] _GEN_86 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],_GEN_74};
  wire  _GEN_87 = RW0_wmask[1];
  wire [43:0] _GEN_88 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    _GEN_74};
  wire  _GEN_89 = RW0_wmask[1];
  wire [44:0] _GEN_90 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],_GEN_74};
  wire [45:0] _GEN_91 = {RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],RW0_wmask[1],
    RW0_wmask[1],RW0_wmask[1],_GEN_74};
  wire  _GEN_92 = ~RW0_wmode;
  wire  _GEN_93 = RW0_wmask[2];
  wire  _GEN_94 = RW0_wmask[2];
  wire  _GEN_95 = RW0_wmask[2];
  wire [1:0] _GEN_96 = {RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_97 = RW0_wmask[2];
  wire [2:0] _GEN_98 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_99 = RW0_wmask[2];
  wire [3:0] _GEN_100 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_101 = RW0_wmask[2];
  wire [4:0] _GEN_102 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_103 = RW0_wmask[2];
  wire [5:0] _GEN_104 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_105 = RW0_wmask[2];
  wire [6:0] _GEN_106 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_107 = RW0_wmask[2];
  wire [7:0] _GEN_108 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2]};
  wire  _GEN_109 = RW0_wmask[2];
  wire [8:0] _GEN_110 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_111 = RW0_wmask[2];
  wire [9:0] _GEN_112 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],RW0_wmask[2],RW0_wmask[2]};
  wire  _GEN_113 = RW0_wmask[2];
  wire [10:0] _GEN_114 = {RW0_wmask[2],_GEN_112};
  wire  _GEN_115 = RW0_wmask[2];
  wire [11:0] _GEN_116 = {RW0_wmask[2],RW0_wmask[2],_GEN_112};
  wire  _GEN_117 = RW0_wmask[2];
  wire [12:0] _GEN_118 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_112};
  wire  _GEN_119 = RW0_wmask[2];
  wire [13:0] _GEN_120 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_112};
  wire  _GEN_121 = RW0_wmask[2];
  wire [14:0] _GEN_122 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_112};
  wire  _GEN_123 = RW0_wmask[2];
  wire [15:0] _GEN_124 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_112};
  wire  _GEN_125 = RW0_wmask[2];
  wire [16:0] _GEN_126 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    _GEN_112};
  wire  _GEN_127 = RW0_wmask[2];
  wire [17:0] _GEN_128 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],_GEN_112};
  wire  _GEN_129 = RW0_wmask[2];
  wire [18:0] _GEN_130 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],RW0_wmask[2],_GEN_112};
  wire  _GEN_131 = RW0_wmask[2];
  wire [19:0] _GEN_132 = {RW0_wmask[2],_GEN_130};
  wire  _GEN_133 = RW0_wmask[2];
  wire [20:0] _GEN_134 = {RW0_wmask[2],RW0_wmask[2],_GEN_130};
  wire  _GEN_135 = RW0_wmask[2];
  wire [21:0] _GEN_136 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_130};
  wire  _GEN_137 = RW0_wmask[3];
  wire [22:0] _GEN_138 = {RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_130};
  wire  _GEN_139 = RW0_wmask[3];
  wire [23:0] _GEN_140 = {RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_130};
  wire  _GEN_141 = RW0_wmask[3];
  wire [24:0] _GEN_142 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],_GEN_130};
  wire  _GEN_143 = RW0_wmask[3];
  wire [25:0] _GEN_144 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    _GEN_130};
  wire  _GEN_145 = RW0_wmask[3];
  wire [26:0] _GEN_146 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],_GEN_130};
  wire  _GEN_147 = RW0_wmask[3];
  wire [27:0] _GEN_148 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[2],RW0_wmask[2],
    RW0_wmask[2],RW0_wmask[2],_GEN_130};
  wire  _GEN_149 = RW0_wmask[3];
  wire [28:0] _GEN_150 = {RW0_wmask[3],_GEN_148};
  wire  _GEN_151 = RW0_wmask[3];
  wire [29:0] _GEN_152 = {RW0_wmask[3],RW0_wmask[3],_GEN_148};
  wire  _GEN_153 = RW0_wmask[3];
  wire [30:0] _GEN_154 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_148};
  wire  _GEN_155 = RW0_wmask[3];
  wire [31:0] _GEN_156 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_148};
  wire  _GEN_157 = RW0_wmask[3];
  wire [32:0] _GEN_158 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_148};
  wire  _GEN_159 = RW0_wmask[3];
  wire [33:0] _GEN_160 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_148};
  wire  _GEN_161 = RW0_wmask[3];
  wire [34:0] _GEN_162 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    _GEN_148};
  wire  _GEN_163 = RW0_wmask[3];
  wire [35:0] _GEN_164 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],_GEN_148};
  wire  _GEN_165 = RW0_wmask[3];
  wire [36:0] _GEN_166 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],RW0_wmask[3],_GEN_148};
  wire  _GEN_167 = RW0_wmask[3];
  wire [37:0] _GEN_168 = {RW0_wmask[3],_GEN_166};
  wire  _GEN_169 = RW0_wmask[3];
  wire [38:0] _GEN_170 = {RW0_wmask[3],RW0_wmask[3],_GEN_166};
  wire  _GEN_171 = RW0_wmask[3];
  wire [39:0] _GEN_172 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_166};
  wire  _GEN_173 = RW0_wmask[3];
  wire [40:0] _GEN_174 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_166};
  wire  _GEN_175 = RW0_wmask[3];
  wire [41:0] _GEN_176 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_166};
  wire  _GEN_177 = RW0_wmask[3];
  wire [42:0] _GEN_178 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],_GEN_166};
  wire  _GEN_179 = RW0_wmask[3];
  wire [43:0] _GEN_180 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    _GEN_166};
  wire  _GEN_181 = RW0_wmask[3];
  wire [44:0] _GEN_182 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],_GEN_166};
  wire [45:0] _GEN_183 = {RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],RW0_wmask[3],
    RW0_wmask[3],RW0_wmask[3],_GEN_166};
  ip224uhdlp1p11rf_512x46m4b2c1s1_t0r0p0d0a1m1h mem_0_0 (
    .adr(mem_0_0_adr),
    .clk(mem_0_0_clk),
    .din(mem_0_0_din),
    .q(mem_0_0_q),
    .ren(mem_0_0_ren),
    .wen(mem_0_0_wen),
    .wbeb(mem_0_0_wbeb),
    .mcen(mem_0_0_mcen),
    .mc(mem_0_0_mc),
    .wa(mem_0_0_wa),
    .wpulse(mem_0_0_wpulse),
    .wpulseen(mem_0_0_wpulseen),
    .fwen(mem_0_0_fwen),
    .clkbyp(mem_0_0_clkbyp)
  );
  ip224uhdlp1p11rf_512x46m4b2c1s1_t0r0p0d0a1m1h mem_0_1 (
    .adr(mem_0_1_adr),
    .clk(mem_0_1_clk),
    .din(mem_0_1_din),
    .q(mem_0_1_q),
    .ren(mem_0_1_ren),
    .wen(mem_0_1_wen),
    .wbeb(mem_0_1_wbeb),
    .mcen(mem_0_1_mcen),
    .mc(mem_0_1_mc),
    .wa(mem_0_1_wa),
    .wpulse(mem_0_1_wpulse),
    .wpulseen(mem_0_1_wpulseen),
    .fwen(mem_0_1_fwen),
    .clkbyp(mem_0_1_clkbyp)
  );
  assign RW0_rdata = {RW0_rdata_0_1,RW0_rdata_0_0};
  assign mem_0_0_adr = {{3'd0}, RW0_addr};
  assign mem_0_0_clk = RW0_clk;
  assign mem_0_0_din = RW0_wdata[45:0];
  assign mem_0_0_ren = ~RW0_wmode & RW0_en;
  assign mem_0_0_wen = RW0_wmode & RW0_en;
  assign mem_0_0_wbeb = ~_GEN_91;
  assign mem_0_0_mcen = 1'h0;
  assign mem_0_0_mc = 3'h0;
  assign mem_0_0_wa = 2'h0;
  assign mem_0_0_wpulse = 2'h0;
  assign mem_0_0_wpulseen = 1'h1;
  assign mem_0_0_fwen = 1'h0;
  assign mem_0_0_clkbyp = 1'h0;
  assign mem_0_1_adr = {{3'd0}, RW0_addr};
  assign mem_0_1_clk = RW0_clk;
  assign mem_0_1_din = RW0_wdata[91:46];
  assign mem_0_1_ren = ~RW0_wmode & RW0_en;
  assign mem_0_1_wen = RW0_wmode & RW0_en;
  assign mem_0_1_wbeb = ~_GEN_183;
  assign mem_0_1_mcen = 1'h0;
  assign mem_0_1_mc = 3'h0;
  assign mem_0_1_wa = 2'h0;
  assign mem_0_1_wpulse = 2'h0;
  assign mem_0_1_wpulseen = 1'h1;
  assign mem_0_1_fwen = 1'h0;
  assign mem_0_1_clkbyp = 1'h0;
endmodule
module dataArrayWay_0_ext(
  input  [8:0]  RW0_addr,
  input         RW0_clk,
  input  [63:0] RW0_wdata,
  output [63:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode
);
  wire [8:0] mem_0_0_adr;
  wire  mem_0_0_clk;
  wire [63:0] mem_0_0_din;
  wire [63:0] mem_0_0_q;
  wire  mem_0_0_ren;
  wire  mem_0_0_wen;
  wire  mem_0_0_mcen;
  wire [2:0] mem_0_0_mc;
  wire [1:0] mem_0_0_wa;
  wire [1:0] mem_0_0_wpulse;
  wire  mem_0_0_wpulseen;
  wire  mem_0_0_fwen;
  wire  mem_0_0_clkbyp;
  wire [63:0] RW0_rdata_0_0 = mem_0_0_q;
  wire [63:0] RW0_rdata_0 = RW0_rdata_0_0;
  wire  _GEN_0 = ~RW0_wmode;
  ip224uhdlp1p11rf_512x64m4b2c1s0_t0r0p0d0a1m1h mem_0_0 (
    .adr(mem_0_0_adr),
    .clk(mem_0_0_clk),
    .din(mem_0_0_din),
    .q(mem_0_0_q),
    .ren(mem_0_0_ren),
    .wen(mem_0_0_wen),
    .mcen(mem_0_0_mcen),
    .mc(mem_0_0_mc),
    .wa(mem_0_0_wa),
    .wpulse(mem_0_0_wpulse),
    .wpulseen(mem_0_0_wpulseen),
    .fwen(mem_0_0_fwen),
    .clkbyp(mem_0_0_clkbyp)
  );
  assign RW0_rdata = mem_0_0_q;
  assign mem_0_0_adr = RW0_addr;
  assign mem_0_0_clk = RW0_clk;
  assign mem_0_0_din = RW0_wdata;
  assign mem_0_0_ren = ~RW0_wmode & RW0_en;
  assign mem_0_0_wen = RW0_wmode & RW0_en;
  assign mem_0_0_mcen = 1'h0;
  assign mem_0_0_mc = 3'h0;
  assign mem_0_0_wa = 2'h0;
  assign mem_0_0_wpulse = 2'h0;
  assign mem_0_0_wpulseen = 1'h1;
  assign mem_0_0_fwen = 1'h0;
  assign mem_0_0_clkbyp = 1'h0;
endmodule
module hi_us_ext(
  input  [7:0] R0_addr,
  input        R0_clk,
  output [3:0] R0_data,
  input        R0_en,
  input  [7:0] W0_addr,
  input        W0_clk,
  input  [3:0] W0_data,
  input        W0_en,
  input  [3:0] W0_mask
);
  wire [7:0] mem_0_0_iarp0;
  wire  mem_0_0_ickrp0;
  wire [3:0] mem_0_0_odoutp0;
  wire  mem_0_0_irenp0;
  wire [7:0] mem_0_0_iawp0;
  wire  mem_0_0_ickwp0;
  wire [3:0] mem_0_0_idinp0;
  wire  mem_0_0_iwenp0;
  wire [3:0] mem_0_0_ibwep0;
  wire  mem_0_0_ifuse;
  wire  mem_0_0_iclkbyp;
  wire  mem_0_0_imce;
  wire [1:0] mem_0_0_irmce;
  wire [3:0] mem_0_0_iwmce;
  wire [3:0] R0_data_0_0 = mem_0_0_odoutp0;
  wire [3:0] R0_data_0 = R0_data_0_0;
  wire  _GEN_0 = W0_mask[1];
  wire  _GEN_1 = W0_mask[0];
  wire  _GEN_2 = W0_mask[2];
  wire [1:0] _GEN_3 = {W0_mask[1],W0_mask[0]};
  wire  _GEN_4 = W0_mask[3];
  wire [2:0] _GEN_5 = {W0_mask[2],W0_mask[1],W0_mask[0]};
  ip224rfsbhpm1r1w256x4be4m1 mem_0_0 (
    .iarp0(mem_0_0_iarp0),
    .ickrp0(mem_0_0_ickrp0),
    .odoutp0(mem_0_0_odoutp0),
    .irenp0(mem_0_0_irenp0),
    .iawp0(mem_0_0_iawp0),
    .ickwp0(mem_0_0_ickwp0),
    .idinp0(mem_0_0_idinp0),
    .iwenp0(mem_0_0_iwenp0),
    .ibwep0(mem_0_0_ibwep0),
    .ifuse(mem_0_0_ifuse),
    .iclkbyp(mem_0_0_iclkbyp),
    .imce(mem_0_0_imce),
    .irmce(mem_0_0_irmce),
    .iwmce(mem_0_0_iwmce)
  );
  assign R0_data = mem_0_0_odoutp0;
  assign mem_0_0_iarp0 = R0_addr;
  assign mem_0_0_ickrp0 = R0_clk;
  assign mem_0_0_irenp0 = R0_en;
  assign mem_0_0_iawp0 = W0_addr;
  assign mem_0_0_ickwp0 = W0_clk;
  assign mem_0_0_idinp0 = W0_data;
  assign mem_0_0_iwenp0 = W0_en;
  assign mem_0_0_ibwep0 = {W0_mask[3],_GEN_5};
  assign mem_0_0_ifuse = 1'h0;
  assign mem_0_0_iclkbyp = 1'h0;
  assign mem_0_0_imce = 1'h0;
  assign mem_0_0_irmce = 2'h0;
  assign mem_0_0_iwmce = 4'h0;
endmodule
module table_ext(
  input  [7:0]  R0_addr,
  input         R0_clk,
  output [43:0] R0_data,
  input         R0_en,
  input  [7:0]  W0_addr,
  input         W0_clk,
  input  [43:0] W0_data,
  input         W0_en,
  input  [3:0]  W0_mask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] mem_0_0_iarp0;
  wire  mem_0_0_ickrp0;
  wire [43:0] mem_0_0_odoutp0;
  wire  mem_0_0_irenp0;
  wire [6:0] mem_0_0_iawp0;
  wire  mem_0_0_ickwp0;
  wire [43:0] mem_0_0_idinp0;
  wire  mem_0_0_iwenp0;
  wire [43:0] mem_0_0_ibwep0;
  wire  mem_0_0_ifuse;
  wire  mem_0_0_iclkbyp;
  wire  mem_0_0_imce;
  wire [1:0] mem_0_0_irmce;
  wire [3:0] mem_0_0_iwmce;
  wire [6:0] mem_1_0_iarp0;
  wire  mem_1_0_ickrp0;
  wire [43:0] mem_1_0_odoutp0;
  wire  mem_1_0_irenp0;
  wire [6:0] mem_1_0_iawp0;
  wire  mem_1_0_ickwp0;
  wire [43:0] mem_1_0_idinp0;
  wire  mem_1_0_iwenp0;
  wire [43:0] mem_1_0_ibwep0;
  wire  mem_1_0_ifuse;
  wire  mem_1_0_iclkbyp;
  wire  mem_1_0_imce;
  wire [1:0] mem_1_0_irmce;
  wire [3:0] mem_1_0_iwmce;
  wire  R0_addr_sel = R0_addr[7];
  reg  R0_addr_sel_reg;
  wire  W0_addr_sel = W0_addr[7];
  wire [43:0] R0_data_0_0 = mem_0_0_odoutp0;
  wire [43:0] R0_data_0 = R0_data_0_0;
  wire [43:0] R0_data_1_0 = mem_1_0_odoutp0;
  wire [43:0] R0_data_1 = R0_data_1_0;
  wire  _GEN_0 = ~R0_addr_sel;
  wire  _GEN_1 = ~W0_addr_sel;
  wire  _GEN_2 = W0_mask[0];
  wire  _GEN_3 = W0_mask[0];
  wire  _GEN_4 = W0_mask[0];
  wire [1:0] _GEN_5 = {W0_mask[0],W0_mask[0]};
  wire  _GEN_6 = W0_mask[0];
  wire [2:0] _GEN_7 = {W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_8 = W0_mask[0];
  wire [3:0] _GEN_9 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_10 = W0_mask[0];
  wire [4:0] _GEN_11 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_12 = W0_mask[0];
  wire [5:0] _GEN_13 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_14 = W0_mask[0];
  wire [6:0] _GEN_15 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_16 = W0_mask[0];
  wire [7:0] _GEN_17 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_18 = W0_mask[0];
  wire [8:0] _GEN_19 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[
    0]};
  wire  _GEN_20 = W0_mask[0];
  wire [9:0] _GEN_21 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[
    0],W0_mask[0]};
  wire  _GEN_22 = W0_mask[1];
  wire [10:0] _GEN_23 = {W0_mask[0],_GEN_21};
  wire  _GEN_24 = W0_mask[1];
  wire [11:0] _GEN_25 = {W0_mask[1],W0_mask[0],_GEN_21};
  wire  _GEN_26 = W0_mask[1];
  wire [12:0] _GEN_27 = {W0_mask[1],W0_mask[1],W0_mask[0],_GEN_21};
  wire  _GEN_28 = W0_mask[1];
  wire [13:0] _GEN_29 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],_GEN_21};
  wire  _GEN_30 = W0_mask[1];
  wire [14:0] _GEN_31 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],_GEN_21};
  wire  _GEN_32 = W0_mask[1];
  wire [15:0] _GEN_33 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],_GEN_21};
  wire  _GEN_34 = W0_mask[1];
  wire [16:0] _GEN_35 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],_GEN_21};
  wire  _GEN_36 = W0_mask[1];
  wire [17:0] _GEN_37 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],_GEN_21
    };
  wire  _GEN_38 = W0_mask[1];
  wire [18:0] _GEN_39 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask
    [0],_GEN_21};
  wire  _GEN_40 = W0_mask[1];
  wire [19:0] _GEN_41 = {W0_mask[1],_GEN_39};
  wire  _GEN_42 = W0_mask[1];
  wire [20:0] _GEN_43 = {W0_mask[1],W0_mask[1],_GEN_39};
  wire  _GEN_44 = W0_mask[2];
  wire [21:0] _GEN_45 = {W0_mask[1],W0_mask[1],W0_mask[1],_GEN_39};
  wire  _GEN_46 = W0_mask[2];
  wire [22:0] _GEN_47 = {W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_39};
  wire  _GEN_48 = W0_mask[2];
  wire [23:0] _GEN_49 = {W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_39};
  wire  _GEN_50 = W0_mask[2];
  wire [24:0] _GEN_51 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_39};
  wire  _GEN_52 = W0_mask[2];
  wire [25:0] _GEN_53 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_39};
  wire  _GEN_54 = W0_mask[2];
  wire [26:0] _GEN_55 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_39
    };
  wire  _GEN_56 = W0_mask[2];
  wire [27:0] _GEN_57 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask
    [1],_GEN_39};
  wire  _GEN_58 = W0_mask[2];
  wire [28:0] _GEN_59 = {W0_mask[2],_GEN_57};
  wire  _GEN_60 = W0_mask[2];
  wire [29:0] _GEN_61 = {W0_mask[2],W0_mask[2],_GEN_57};
  wire  _GEN_62 = W0_mask[2];
  wire [30:0] _GEN_63 = {W0_mask[2],W0_mask[2],W0_mask[2],_GEN_57};
  wire  _GEN_64 = W0_mask[2];
  wire [31:0] _GEN_65 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_57};
  wire  _GEN_66 = W0_mask[3];
  wire [32:0] _GEN_67 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_57};
  wire  _GEN_68 = W0_mask[3];
  wire [33:0] _GEN_69 = {W0_mask[3],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_57};
  wire  _GEN_70 = W0_mask[3];
  wire [34:0] _GEN_71 = {W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_57};
  wire  _GEN_72 = W0_mask[3];
  wire [35:0] _GEN_73 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_57
    };
  wire  _GEN_74 = W0_mask[3];
  wire [36:0] _GEN_75 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask
    [2],_GEN_57};
  wire  _GEN_76 = W0_mask[3];
  wire [37:0] _GEN_77 = {W0_mask[3],_GEN_75};
  wire  _GEN_78 = W0_mask[3];
  wire [38:0] _GEN_79 = {W0_mask[3],W0_mask[3],_GEN_75};
  wire  _GEN_80 = W0_mask[3];
  wire [39:0] _GEN_81 = {W0_mask[3],W0_mask[3],W0_mask[3],_GEN_75};
  wire  _GEN_82 = W0_mask[3];
  wire [40:0] _GEN_83 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_75};
  wire  _GEN_84 = W0_mask[3];
  wire [41:0] _GEN_85 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_75};
  wire  _GEN_86 = W0_mask[3];
  wire [42:0] _GEN_87 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_75};
  wire  _GEN_88 = W0_mask[0];
  wire  _GEN_89 = W0_mask[0];
  wire  _GEN_90 = W0_mask[0];
  wire [1:0] _GEN_91 = {W0_mask[0],W0_mask[0]};
  wire  _GEN_92 = W0_mask[0];
  wire [2:0] _GEN_93 = {W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_94 = W0_mask[0];
  wire [3:0] _GEN_95 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_96 = W0_mask[0];
  wire [4:0] _GEN_97 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_98 = W0_mask[0];
  wire [5:0] _GEN_99 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_100 = W0_mask[0];
  wire [6:0] _GEN_101 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_102 = W0_mask[0];
  wire [7:0] _GEN_103 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_104 = W0_mask[0];
  wire [8:0] _GEN_105 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask
    [0]};
  wire  _GEN_106 = W0_mask[0];
  wire [9:0] _GEN_107 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask
    [0],W0_mask[0]};
  wire  _GEN_108 = W0_mask[1];
  wire [10:0] _GEN_109 = {W0_mask[0],_GEN_21};
  wire  _GEN_110 = W0_mask[1];
  wire [11:0] _GEN_111 = {W0_mask[1],W0_mask[0],_GEN_21};
  wire  _GEN_112 = W0_mask[1];
  wire [12:0] _GEN_113 = {W0_mask[1],W0_mask[1],W0_mask[0],_GEN_21};
  wire  _GEN_114 = W0_mask[1];
  wire [13:0] _GEN_115 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],_GEN_21};
  wire  _GEN_116 = W0_mask[1];
  wire [14:0] _GEN_117 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],_GEN_21};
  wire  _GEN_118 = W0_mask[1];
  wire [15:0] _GEN_119 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],_GEN_21};
  wire  _GEN_120 = W0_mask[1];
  wire [16:0] _GEN_121 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],_GEN_21};
  wire  _GEN_122 = W0_mask[1];
  wire [17:0] _GEN_123 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],
    _GEN_21};
  wire  _GEN_124 = W0_mask[1];
  wire [18:0] _GEN_125 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],
    W0_mask[0],_GEN_21};
  wire  _GEN_126 = W0_mask[1];
  wire [19:0] _GEN_127 = {W0_mask[1],_GEN_39};
  wire  _GEN_128 = W0_mask[1];
  wire [20:0] _GEN_129 = {W0_mask[1],W0_mask[1],_GEN_39};
  wire  _GEN_130 = W0_mask[2];
  wire [21:0] _GEN_131 = {W0_mask[1],W0_mask[1],W0_mask[1],_GEN_39};
  wire  _GEN_132 = W0_mask[2];
  wire [22:0] _GEN_133 = {W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_39};
  wire  _GEN_134 = W0_mask[2];
  wire [23:0] _GEN_135 = {W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_39};
  wire  _GEN_136 = W0_mask[2];
  wire [24:0] _GEN_137 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_39};
  wire  _GEN_138 = W0_mask[2];
  wire [25:0] _GEN_139 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_39};
  wire  _GEN_140 = W0_mask[2];
  wire [26:0] _GEN_141 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],
    _GEN_39};
  wire  _GEN_142 = W0_mask[2];
  wire [27:0] _GEN_143 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],
    W0_mask[1],_GEN_39};
  wire  _GEN_144 = W0_mask[2];
  wire [28:0] _GEN_145 = {W0_mask[2],_GEN_57};
  wire  _GEN_146 = W0_mask[2];
  wire [29:0] _GEN_147 = {W0_mask[2],W0_mask[2],_GEN_57};
  wire  _GEN_148 = W0_mask[2];
  wire [30:0] _GEN_149 = {W0_mask[2],W0_mask[2],W0_mask[2],_GEN_57};
  wire  _GEN_150 = W0_mask[2];
  wire [31:0] _GEN_151 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_57};
  wire  _GEN_152 = W0_mask[3];
  wire [32:0] _GEN_153 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_57};
  wire  _GEN_154 = W0_mask[3];
  wire [33:0] _GEN_155 = {W0_mask[3],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_57};
  wire  _GEN_156 = W0_mask[3];
  wire [34:0] _GEN_157 = {W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_57};
  wire  _GEN_158 = W0_mask[3];
  wire [35:0] _GEN_159 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],
    _GEN_57};
  wire  _GEN_160 = W0_mask[3];
  wire [36:0] _GEN_161 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],
    W0_mask[2],_GEN_57};
  wire  _GEN_162 = W0_mask[3];
  wire [37:0] _GEN_163 = {W0_mask[3],_GEN_75};
  wire  _GEN_164 = W0_mask[3];
  wire [38:0] _GEN_165 = {W0_mask[3],W0_mask[3],_GEN_75};
  wire  _GEN_166 = W0_mask[3];
  wire [39:0] _GEN_167 = {W0_mask[3],W0_mask[3],W0_mask[3],_GEN_75};
  wire  _GEN_168 = W0_mask[3];
  wire [40:0] _GEN_169 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_75};
  wire  _GEN_170 = W0_mask[3];
  wire [41:0] _GEN_171 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_75};
  wire  _GEN_172 = W0_mask[3];
  wire [42:0] _GEN_173 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_75};
  ip224rfsbhpm1r1w128x44be44m1 mem_0_0 (
    .iarp0(mem_0_0_iarp0),
    .ickrp0(mem_0_0_ickrp0),
    .odoutp0(mem_0_0_odoutp0),
    .irenp0(mem_0_0_irenp0),
    .iawp0(mem_0_0_iawp0),
    .ickwp0(mem_0_0_ickwp0),
    .idinp0(mem_0_0_idinp0),
    .iwenp0(mem_0_0_iwenp0),
    .ibwep0(mem_0_0_ibwep0),
    .ifuse(mem_0_0_ifuse),
    .iclkbyp(mem_0_0_iclkbyp),
    .imce(mem_0_0_imce),
    .irmce(mem_0_0_irmce),
    .iwmce(mem_0_0_iwmce)
  );
  ip224rfsbhpm1r1w128x44be44m1 mem_1_0 (
    .iarp0(mem_1_0_iarp0),
    .ickrp0(mem_1_0_ickrp0),
    .odoutp0(mem_1_0_odoutp0),
    .irenp0(mem_1_0_irenp0),
    .iawp0(mem_1_0_iawp0),
    .ickwp0(mem_1_0_ickwp0),
    .idinp0(mem_1_0_idinp0),
    .iwenp0(mem_1_0_iwenp0),
    .ibwep0(mem_1_0_ibwep0),
    .ifuse(mem_1_0_ifuse),
    .iclkbyp(mem_1_0_iclkbyp),
    .imce(mem_1_0_imce),
    .irmce(mem_1_0_irmce),
    .iwmce(mem_1_0_iwmce)
  );
  assign R0_data = ~R0_addr_sel_reg ? R0_data_0_0 : R0_addr_sel_reg ? R0_data_1_0 : 44'h0;
  assign mem_0_0_iarp0 = R0_addr[6:0];
  assign mem_0_0_ickrp0 = R0_clk;
  assign mem_0_0_irenp0 = R0_en & ~R0_addr_sel;
  assign mem_0_0_iawp0 = W0_addr[6:0];
  assign mem_0_0_ickwp0 = W0_clk;
  assign mem_0_0_idinp0 = W0_data;
  assign mem_0_0_iwenp0 = W0_en & ~W0_addr_sel;
  assign mem_0_0_ibwep0 = {W0_mask[3],_GEN_87};
  assign mem_0_0_ifuse = 1'h0;
  assign mem_0_0_iclkbyp = 1'h0;
  assign mem_0_0_imce = 1'h0;
  assign mem_0_0_irmce = 2'h0;
  assign mem_0_0_iwmce = 4'h0;
  assign mem_1_0_iarp0 = R0_addr[6:0];
  assign mem_1_0_ickrp0 = R0_clk;
  assign mem_1_0_irenp0 = R0_en & R0_addr_sel;
  assign mem_1_0_iawp0 = W0_addr[6:0];
  assign mem_1_0_ickwp0 = W0_clk;
  assign mem_1_0_idinp0 = W0_data;
  assign mem_1_0_iwenp0 = W0_en & W0_addr_sel;
  assign mem_1_0_ibwep0 = {W0_mask[3],_GEN_87};
  assign mem_1_0_ifuse = 1'h0;
  assign mem_1_0_iclkbyp = 1'h0;
  assign mem_1_0_imce = 1'h0;
  assign mem_1_0_irmce = 2'h0;
  assign mem_1_0_iwmce = 4'h0;
  always @(posedge R0_clk) begin
    if (R0_en) begin
      R0_addr_sel_reg <= R0_addr_sel;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  R0_addr_sel_reg = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module meta_0_ext(
  input  [6:0]   R0_addr,
  input          R0_clk,
  output [123:0] R0_data,
  input          R0_en,
  input  [6:0]   W0_addr,
  input          W0_clk,
  input  [123:0] W0_data,
  input          W0_en,
  input  [3:0]   W0_mask
);
  wire [6:0] mem_0_0_iarp0;
  wire  mem_0_0_ickrp0;
  wire [123:0] mem_0_0_odoutp0;
  wire  mem_0_0_irenp0;
  wire [6:0] mem_0_0_iawp0;
  wire  mem_0_0_ickwp0;
  wire [123:0] mem_0_0_idinp0;
  wire  mem_0_0_iwenp0;
  wire [123:0] mem_0_0_ibwep0;
  wire  mem_0_0_ifuse;
  wire  mem_0_0_iclkbyp;
  wire  mem_0_0_imce;
  wire [1:0] mem_0_0_irmce;
  wire [3:0] mem_0_0_iwmce;
  wire [123:0] R0_data_0_0 = mem_0_0_odoutp0;
  wire [123:0] R0_data_0 = R0_data_0_0;
  wire  _GEN_0 = W0_mask[0];
  wire  _GEN_1 = W0_mask[0];
  wire  _GEN_2 = W0_mask[0];
  wire [1:0] _GEN_3 = {W0_mask[0],W0_mask[0]};
  wire  _GEN_4 = W0_mask[0];
  wire [2:0] _GEN_5 = {W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_6 = W0_mask[0];
  wire [3:0] _GEN_7 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_8 = W0_mask[0];
  wire [4:0] _GEN_9 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_10 = W0_mask[0];
  wire [5:0] _GEN_11 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_12 = W0_mask[0];
  wire [6:0] _GEN_13 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_14 = W0_mask[0];
  wire [7:0] _GEN_15 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_16 = W0_mask[0];
  wire [8:0] _GEN_17 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[
    0]};
  wire  _GEN_18 = W0_mask[0];
  wire [9:0] _GEN_19 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[
    0],W0_mask[0]};
  wire  _GEN_20 = W0_mask[0];
  wire [10:0] _GEN_21 = {W0_mask[0],_GEN_19};
  wire  _GEN_22 = W0_mask[0];
  wire [11:0] _GEN_23 = {W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_24 = W0_mask[0];
  wire [12:0] _GEN_25 = {W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_26 = W0_mask[0];
  wire [13:0] _GEN_27 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_28 = W0_mask[0];
  wire [14:0] _GEN_29 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_30 = W0_mask[0];
  wire [15:0] _GEN_31 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_32 = W0_mask[0];
  wire [16:0] _GEN_33 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_34 = W0_mask[0];
  wire [17:0] _GEN_35 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19
    };
  wire  _GEN_36 = W0_mask[0];
  wire [18:0] _GEN_37 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask
    [0],_GEN_19};
  wire  _GEN_38 = W0_mask[0];
  wire [19:0] _GEN_39 = {W0_mask[0],_GEN_37};
  wire  _GEN_40 = W0_mask[0];
  wire [20:0] _GEN_41 = {W0_mask[0],W0_mask[0],_GEN_37};
  wire  _GEN_42 = W0_mask[0];
  wire [21:0] _GEN_43 = {W0_mask[0],W0_mask[0],W0_mask[0],_GEN_37};
  wire  _GEN_44 = W0_mask[0];
  wire [22:0] _GEN_45 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_37};
  wire  _GEN_46 = W0_mask[0];
  wire [23:0] _GEN_47 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_37};
  wire  _GEN_48 = W0_mask[0];
  wire [24:0] _GEN_49 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_37};
  wire  _GEN_50 = W0_mask[0];
  wire [25:0] _GEN_51 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_37};
  wire  _GEN_52 = W0_mask[0];
  wire [26:0] _GEN_53 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_37
    };
  wire  _GEN_54 = W0_mask[0];
  wire [27:0] _GEN_55 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask
    [0],_GEN_37};
  wire  _GEN_56 = W0_mask[0];
  wire [28:0] _GEN_57 = {W0_mask[0],_GEN_55};
  wire  _GEN_58 = W0_mask[0];
  wire [29:0] _GEN_59 = {W0_mask[0],W0_mask[0],_GEN_55};
  wire  _GEN_60 = W0_mask[1];
  wire [30:0] _GEN_61 = {W0_mask[0],W0_mask[0],W0_mask[0],_GEN_55};
  wire  _GEN_62 = W0_mask[1];
  wire [31:0] _GEN_63 = {W0_mask[1],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_55};
  wire  _GEN_64 = W0_mask[1];
  wire [32:0] _GEN_65 = {W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_55};
  wire  _GEN_66 = W0_mask[1];
  wire [33:0] _GEN_67 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_55};
  wire  _GEN_68 = W0_mask[1];
  wire [34:0] _GEN_69 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_55};
  wire  _GEN_70 = W0_mask[1];
  wire [35:0] _GEN_71 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_55
    };
  wire  _GEN_72 = W0_mask[1];
  wire [36:0] _GEN_73 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0],W0_mask
    [0],_GEN_55};
  wire  _GEN_74 = W0_mask[1];
  wire [37:0] _GEN_75 = {W0_mask[1],_GEN_73};
  wire  _GEN_76 = W0_mask[1];
  wire [38:0] _GEN_77 = {W0_mask[1],W0_mask[1],_GEN_73};
  wire  _GEN_78 = W0_mask[1];
  wire [39:0] _GEN_79 = {W0_mask[1],W0_mask[1],W0_mask[1],_GEN_73};
  wire  _GEN_80 = W0_mask[1];
  wire [40:0] _GEN_81 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_73};
  wire  _GEN_82 = W0_mask[1];
  wire [41:0] _GEN_83 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_73};
  wire  _GEN_84 = W0_mask[1];
  wire [42:0] _GEN_85 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_73};
  wire  _GEN_86 = W0_mask[1];
  wire [43:0] _GEN_87 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_73};
  wire  _GEN_88 = W0_mask[1];
  wire [44:0] _GEN_89 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_73
    };
  wire  _GEN_90 = W0_mask[1];
  wire [45:0] _GEN_91 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask
    [1],_GEN_73};
  wire  _GEN_92 = W0_mask[1];
  wire [46:0] _GEN_93 = {W0_mask[1],_GEN_91};
  wire  _GEN_94 = W0_mask[1];
  wire [47:0] _GEN_95 = {W0_mask[1],W0_mask[1],_GEN_91};
  wire  _GEN_96 = W0_mask[1];
  wire [48:0] _GEN_97 = {W0_mask[1],W0_mask[1],W0_mask[1],_GEN_91};
  wire  _GEN_98 = W0_mask[1];
  wire [49:0] _GEN_99 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_91};
  wire  _GEN_100 = W0_mask[1];
  wire [50:0] _GEN_101 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_91};
  wire  _GEN_102 = W0_mask[1];
  wire [51:0] _GEN_103 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_91};
  wire  _GEN_104 = W0_mask[1];
  wire [52:0] _GEN_105 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_91};
  wire  _GEN_106 = W0_mask[1];
  wire [53:0] _GEN_107 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],
    _GEN_91};
  wire  _GEN_108 = W0_mask[1];
  wire [54:0] _GEN_109 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],
    W0_mask[1],_GEN_91};
  wire  _GEN_110 = W0_mask[1];
  wire [55:0] _GEN_111 = {W0_mask[1],_GEN_109};
  wire  _GEN_112 = W0_mask[1];
  wire [56:0] _GEN_113 = {W0_mask[1],W0_mask[1],_GEN_109};
  wire  _GEN_114 = W0_mask[1];
  wire [57:0] _GEN_115 = {W0_mask[1],W0_mask[1],W0_mask[1],_GEN_109};
  wire  _GEN_116 = W0_mask[1];
  wire [58:0] _GEN_117 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_109};
  wire  _GEN_118 = W0_mask[1];
  wire [59:0] _GEN_119 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_109};
  wire  _GEN_120 = W0_mask[1];
  wire [60:0] _GEN_121 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_109};
  wire  _GEN_122 = W0_mask[2];
  wire [61:0] _GEN_123 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_109};
  wire  _GEN_124 = W0_mask[2];
  wire [62:0] _GEN_125 = {W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],
    _GEN_109};
  wire  _GEN_126 = W0_mask[2];
  wire [63:0] _GEN_127 = {W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],
    W0_mask[1],_GEN_109};
  wire  _GEN_128 = W0_mask[2];
  wire [64:0] _GEN_129 = {W0_mask[2],_GEN_127};
  wire  _GEN_130 = W0_mask[2];
  wire [65:0] _GEN_131 = {W0_mask[2],W0_mask[2],_GEN_127};
  wire  _GEN_132 = W0_mask[2];
  wire [66:0] _GEN_133 = {W0_mask[2],W0_mask[2],W0_mask[2],_GEN_127};
  wire  _GEN_134 = W0_mask[2];
  wire [67:0] _GEN_135 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_127};
  wire  _GEN_136 = W0_mask[2];
  wire [68:0] _GEN_137 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_127};
  wire  _GEN_138 = W0_mask[2];
  wire [69:0] _GEN_139 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_127};
  wire  _GEN_140 = W0_mask[2];
  wire [70:0] _GEN_141 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_127};
  wire  _GEN_142 = W0_mask[2];
  wire [71:0] _GEN_143 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],
    _GEN_127};
  wire  _GEN_144 = W0_mask[2];
  wire [72:0] _GEN_145 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],
    W0_mask[2],_GEN_127};
  wire  _GEN_146 = W0_mask[2];
  wire [73:0] _GEN_147 = {W0_mask[2],_GEN_145};
  wire  _GEN_148 = W0_mask[2];
  wire [74:0] _GEN_149 = {W0_mask[2],W0_mask[2],_GEN_145};
  wire  _GEN_150 = W0_mask[2];
  wire [75:0] _GEN_151 = {W0_mask[2],W0_mask[2],W0_mask[2],_GEN_145};
  wire  _GEN_152 = W0_mask[2];
  wire [76:0] _GEN_153 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_145};
  wire  _GEN_154 = W0_mask[2];
  wire [77:0] _GEN_155 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_145};
  wire  _GEN_156 = W0_mask[2];
  wire [78:0] _GEN_157 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_145};
  wire  _GEN_158 = W0_mask[2];
  wire [79:0] _GEN_159 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_145};
  wire  _GEN_160 = W0_mask[2];
  wire [80:0] _GEN_161 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],
    _GEN_145};
  wire  _GEN_162 = W0_mask[2];
  wire [81:0] _GEN_163 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],
    W0_mask[2],_GEN_145};
  wire  _GEN_164 = W0_mask[2];
  wire [82:0] _GEN_165 = {W0_mask[2],_GEN_163};
  wire  _GEN_166 = W0_mask[2];
  wire [83:0] _GEN_167 = {W0_mask[2],W0_mask[2],_GEN_163};
  wire  _GEN_168 = W0_mask[2];
  wire [84:0] _GEN_169 = {W0_mask[2],W0_mask[2],W0_mask[2],_GEN_163};
  wire  _GEN_170 = W0_mask[2];
  wire [85:0] _GEN_171 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_163};
  wire  _GEN_172 = W0_mask[2];
  wire [86:0] _GEN_173 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_163};
  wire  _GEN_174 = W0_mask[2];
  wire [87:0] _GEN_175 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_163};
  wire  _GEN_176 = W0_mask[2];
  wire [88:0] _GEN_177 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_163};
  wire  _GEN_178 = W0_mask[2];
  wire [89:0] _GEN_179 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],
    _GEN_163};
  wire  _GEN_180 = W0_mask[2];
  wire [90:0] _GEN_181 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],
    W0_mask[2],_GEN_163};
  wire  _GEN_182 = W0_mask[2];
  wire [91:0] _GEN_183 = {W0_mask[2],_GEN_181};
  wire  _GEN_184 = W0_mask[3];
  wire [92:0] _GEN_185 = {W0_mask[2],W0_mask[2],_GEN_181};
  wire  _GEN_186 = W0_mask[3];
  wire [93:0] _GEN_187 = {W0_mask[3],W0_mask[2],W0_mask[2],_GEN_181};
  wire  _GEN_188 = W0_mask[3];
  wire [94:0] _GEN_189 = {W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],_GEN_181};
  wire  _GEN_190 = W0_mask[3];
  wire [95:0] _GEN_191 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],_GEN_181};
  wire  _GEN_192 = W0_mask[3];
  wire [96:0] _GEN_193 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],_GEN_181};
  wire  _GEN_194 = W0_mask[3];
  wire [97:0] _GEN_195 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],_GEN_181};
  wire  _GEN_196 = W0_mask[3];
  wire [98:0] _GEN_197 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],
    _GEN_181};
  wire  _GEN_198 = W0_mask[3];
  wire [99:0] _GEN_199 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],
    W0_mask[2],_GEN_181};
  wire  _GEN_200 = W0_mask[3];
  wire [100:0] _GEN_201 = {W0_mask[3],_GEN_199};
  wire  _GEN_202 = W0_mask[3];
  wire [101:0] _GEN_203 = {W0_mask[3],W0_mask[3],_GEN_199};
  wire  _GEN_204 = W0_mask[3];
  wire [102:0] _GEN_205 = {W0_mask[3],W0_mask[3],W0_mask[3],_GEN_199};
  wire  _GEN_206 = W0_mask[3];
  wire [103:0] _GEN_207 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_199};
  wire  _GEN_208 = W0_mask[3];
  wire [104:0] _GEN_209 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_199};
  wire  _GEN_210 = W0_mask[3];
  wire [105:0] _GEN_211 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_199};
  wire  _GEN_212 = W0_mask[3];
  wire [106:0] _GEN_213 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_199};
  wire  _GEN_214 = W0_mask[3];
  wire [107:0] _GEN_215 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],
    _GEN_199};
  wire  _GEN_216 = W0_mask[3];
  wire [108:0] _GEN_217 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],
    W0_mask[3],_GEN_199};
  wire  _GEN_218 = W0_mask[3];
  wire [109:0] _GEN_219 = {W0_mask[3],_GEN_217};
  wire  _GEN_220 = W0_mask[3];
  wire [110:0] _GEN_221 = {W0_mask[3],W0_mask[3],_GEN_217};
  wire  _GEN_222 = W0_mask[3];
  wire [111:0] _GEN_223 = {W0_mask[3],W0_mask[3],W0_mask[3],_GEN_217};
  wire  _GEN_224 = W0_mask[3];
  wire [112:0] _GEN_225 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_217};
  wire  _GEN_226 = W0_mask[3];
  wire [113:0] _GEN_227 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_217};
  wire  _GEN_228 = W0_mask[3];
  wire [114:0] _GEN_229 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_217};
  wire  _GEN_230 = W0_mask[3];
  wire [115:0] _GEN_231 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_217};
  wire  _GEN_232 = W0_mask[3];
  wire [116:0] _GEN_233 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],
    _GEN_217};
  wire  _GEN_234 = W0_mask[3];
  wire [117:0] _GEN_235 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],
    W0_mask[3],_GEN_217};
  wire  _GEN_236 = W0_mask[3];
  wire [118:0] _GEN_237 = {W0_mask[3],_GEN_235};
  wire  _GEN_238 = W0_mask[3];
  wire [119:0] _GEN_239 = {W0_mask[3],W0_mask[3],_GEN_235};
  wire  _GEN_240 = W0_mask[3];
  wire [120:0] _GEN_241 = {W0_mask[3],W0_mask[3],W0_mask[3],_GEN_235};
  wire  _GEN_242 = W0_mask[3];
  wire [121:0] _GEN_243 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_235};
  wire  _GEN_244 = W0_mask[3];
  wire [122:0] _GEN_245 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_235};
  ip224rfsbhpm1r1w128x124be124m1 mem_0_0 (
    .iarp0(mem_0_0_iarp0),
    .ickrp0(mem_0_0_ickrp0),
    .odoutp0(mem_0_0_odoutp0),
    .irenp0(mem_0_0_irenp0),
    .iawp0(mem_0_0_iawp0),
    .ickwp0(mem_0_0_ickwp0),
    .idinp0(mem_0_0_idinp0),
    .iwenp0(mem_0_0_iwenp0),
    .ibwep0(mem_0_0_ibwep0),
    .ifuse(mem_0_0_ifuse),
    .iclkbyp(mem_0_0_iclkbyp),
    .imce(mem_0_0_imce),
    .irmce(mem_0_0_irmce),
    .iwmce(mem_0_0_iwmce)
  );
  assign R0_data = mem_0_0_odoutp0;
  assign mem_0_0_iarp0 = R0_addr;
  assign mem_0_0_ickrp0 = R0_clk;
  assign mem_0_0_irenp0 = R0_en;
  assign mem_0_0_iawp0 = W0_addr;
  assign mem_0_0_ickwp0 = W0_clk;
  assign mem_0_0_idinp0 = W0_data;
  assign mem_0_0_iwenp0 = W0_en;
  assign mem_0_0_ibwep0 = {W0_mask[3],_GEN_245};
  assign mem_0_0_ifuse = 1'h0;
  assign mem_0_0_iclkbyp = 1'h0;
  assign mem_0_0_imce = 1'h0;
  assign mem_0_0_irmce = 2'h0;
  assign mem_0_0_iwmce = 4'h0;
endmodule
module btb_0_ext(
  input  [6:0]  R0_addr,
  input         R0_clk,
  output [55:0] R0_data,
  input         R0_en,
  input  [6:0]  W0_addr,
  input         W0_clk,
  input  [55:0] W0_data,
  input         W0_en,
  input  [3:0]  W0_mask
);
  wire [6:0] mem_0_0_iarp0;
  wire  mem_0_0_ickrp0;
  wire [55:0] mem_0_0_odoutp0;
  wire  mem_0_0_irenp0;
  wire [6:0] mem_0_0_iawp0;
  wire  mem_0_0_ickwp0;
  wire [55:0] mem_0_0_idinp0;
  wire  mem_0_0_iwenp0;
  wire [55:0] mem_0_0_ibwep0;
  wire  mem_0_0_ifuse;
  wire  mem_0_0_iclkbyp;
  wire  mem_0_0_imce;
  wire [1:0] mem_0_0_irmce;
  wire [3:0] mem_0_0_iwmce;
  wire [55:0] R0_data_0_0 = mem_0_0_odoutp0;
  wire [55:0] R0_data_0 = R0_data_0_0;
  wire  _GEN_0 = W0_mask[0];
  wire  _GEN_1 = W0_mask[0];
  wire  _GEN_2 = W0_mask[0];
  wire [1:0] _GEN_3 = {W0_mask[0],W0_mask[0]};
  wire  _GEN_4 = W0_mask[0];
  wire [2:0] _GEN_5 = {W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_6 = W0_mask[0];
  wire [3:0] _GEN_7 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_8 = W0_mask[0];
  wire [4:0] _GEN_9 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_10 = W0_mask[0];
  wire [5:0] _GEN_11 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_12 = W0_mask[0];
  wire [6:0] _GEN_13 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_14 = W0_mask[0];
  wire [7:0] _GEN_15 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0]};
  wire  _GEN_16 = W0_mask[0];
  wire [8:0] _GEN_17 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[
    0]};
  wire  _GEN_18 = W0_mask[0];
  wire [9:0] _GEN_19 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[
    0],W0_mask[0]};
  wire  _GEN_20 = W0_mask[0];
  wire [10:0] _GEN_21 = {W0_mask[0],_GEN_19};
  wire  _GEN_22 = W0_mask[0];
  wire [11:0] _GEN_23 = {W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_24 = W0_mask[0];
  wire [12:0] _GEN_25 = {W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_26 = W0_mask[1];
  wire [13:0] _GEN_27 = {W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_28 = W0_mask[1];
  wire [14:0] _GEN_29 = {W0_mask[1],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_30 = W0_mask[1];
  wire [15:0] _GEN_31 = {W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_32 = W0_mask[1];
  wire [16:0] _GEN_33 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19};
  wire  _GEN_34 = W0_mask[1];
  wire [17:0] _GEN_35 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask[0],_GEN_19
    };
  wire  _GEN_36 = W0_mask[1];
  wire [18:0] _GEN_37 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0],W0_mask[0],W0_mask
    [0],_GEN_19};
  wire  _GEN_38 = W0_mask[1];
  wire [19:0] _GEN_39 = {W0_mask[1],_GEN_37};
  wire  _GEN_40 = W0_mask[1];
  wire [20:0] _GEN_41 = {W0_mask[1],W0_mask[1],_GEN_37};
  wire  _GEN_42 = W0_mask[1];
  wire [21:0] _GEN_43 = {W0_mask[1],W0_mask[1],W0_mask[1],_GEN_37};
  wire  _GEN_44 = W0_mask[1];
  wire [22:0] _GEN_45 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_37};
  wire  _GEN_46 = W0_mask[1];
  wire [23:0] _GEN_47 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_37};
  wire  _GEN_48 = W0_mask[1];
  wire [24:0] _GEN_49 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_37};
  wire  _GEN_50 = W0_mask[1];
  wire [25:0] _GEN_51 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_37};
  wire  _GEN_52 = W0_mask[1];
  wire [26:0] _GEN_53 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],_GEN_37
    };
  wire  _GEN_54 = W0_mask[2];
  wire [27:0] _GEN_55 = {W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask[1],W0_mask
    [1],_GEN_37};
  wire  _GEN_56 = W0_mask[2];
  wire [28:0] _GEN_57 = {W0_mask[2],_GEN_55};
  wire  _GEN_58 = W0_mask[2];
  wire [29:0] _GEN_59 = {W0_mask[2],W0_mask[2],_GEN_55};
  wire  _GEN_60 = W0_mask[2];
  wire [30:0] _GEN_61 = {W0_mask[2],W0_mask[2],W0_mask[2],_GEN_55};
  wire  _GEN_62 = W0_mask[2];
  wire [31:0] _GEN_63 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_55};
  wire  _GEN_64 = W0_mask[2];
  wire [32:0] _GEN_65 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_55};
  wire  _GEN_66 = W0_mask[2];
  wire [33:0] _GEN_67 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_55};
  wire  _GEN_68 = W0_mask[2];
  wire [34:0] _GEN_69 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_55};
  wire  _GEN_70 = W0_mask[2];
  wire [35:0] _GEN_71 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_55
    };
  wire  _GEN_72 = W0_mask[2];
  wire [36:0] _GEN_73 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask
    [2],_GEN_55};
  wire  _GEN_74 = W0_mask[2];
  wire [37:0] _GEN_75 = {W0_mask[2],_GEN_73};
  wire  _GEN_76 = W0_mask[2];
  wire [38:0] _GEN_77 = {W0_mask[2],W0_mask[2],_GEN_73};
  wire  _GEN_78 = W0_mask[2];
  wire [39:0] _GEN_79 = {W0_mask[2],W0_mask[2],W0_mask[2],_GEN_73};
  wire  _GEN_80 = W0_mask[2];
  wire [40:0] _GEN_81 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_73};
  wire  _GEN_82 = W0_mask[3];
  wire [41:0] _GEN_83 = {W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_73};
  wire  _GEN_84 = W0_mask[3];
  wire [42:0] _GEN_85 = {W0_mask[3],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_73};
  wire  _GEN_86 = W0_mask[3];
  wire [43:0] _GEN_87 = {W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_73};
  wire  _GEN_88 = W0_mask[3];
  wire [44:0] _GEN_89 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],_GEN_73
    };
  wire  _GEN_90 = W0_mask[3];
  wire [45:0] _GEN_91 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask[2],W0_mask
    [2],_GEN_73};
  wire  _GEN_92 = W0_mask[3];
  wire [46:0] _GEN_93 = {W0_mask[3],_GEN_91};
  wire  _GEN_94 = W0_mask[3];
  wire [47:0] _GEN_95 = {W0_mask[3],W0_mask[3],_GEN_91};
  wire  _GEN_96 = W0_mask[3];
  wire [48:0] _GEN_97 = {W0_mask[3],W0_mask[3],W0_mask[3],_GEN_91};
  wire  _GEN_98 = W0_mask[3];
  wire [49:0] _GEN_99 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_91};
  wire  _GEN_100 = W0_mask[3];
  wire [50:0] _GEN_101 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_91};
  wire  _GEN_102 = W0_mask[3];
  wire [51:0] _GEN_103 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_91};
  wire  _GEN_104 = W0_mask[3];
  wire [52:0] _GEN_105 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],_GEN_91};
  wire  _GEN_106 = W0_mask[3];
  wire [53:0] _GEN_107 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],
    _GEN_91};
  wire  _GEN_108 = W0_mask[3];
  wire [54:0] _GEN_109 = {W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],W0_mask[3],
    W0_mask[3],_GEN_91};
  ip224rfsbhpm1r1w128x56be56m1 mem_0_0 (
    .iarp0(mem_0_0_iarp0),
    .ickrp0(mem_0_0_ickrp0),
    .odoutp0(mem_0_0_odoutp0),
    .irenp0(mem_0_0_irenp0),
    .iawp0(mem_0_0_iawp0),
    .ickwp0(mem_0_0_ickwp0),
    .idinp0(mem_0_0_idinp0),
    .iwenp0(mem_0_0_iwenp0),
    .ibwep0(mem_0_0_ibwep0),
    .ifuse(mem_0_0_ifuse),
    .iclkbyp(mem_0_0_iclkbyp),
    .imce(mem_0_0_imce),
    .irmce(mem_0_0_irmce),
    .iwmce(mem_0_0_iwmce)
  );
  assign R0_data = mem_0_0_odoutp0;
  assign mem_0_0_iarp0 = R0_addr;
  assign mem_0_0_ickrp0 = R0_clk;
  assign mem_0_0_irenp0 = R0_en;
  assign mem_0_0_iawp0 = W0_addr;
  assign mem_0_0_ickwp0 = W0_clk;
  assign mem_0_0_idinp0 = W0_data;
  assign mem_0_0_iwenp0 = W0_en;
  assign mem_0_0_ibwep0 = {W0_mask[3],_GEN_109};
  assign mem_0_0_ifuse = 1'h0;
  assign mem_0_0_iclkbyp = 1'h0;
  assign mem_0_0_imce = 1'h0;
  assign mem_0_0_irmce = 2'h0;
  assign mem_0_0_iwmce = 4'h0;
endmodule
module ebtb_ext(
  input  [6:0]  R0_addr,
  input         R0_clk,
  output [39:0] R0_data,
  input         R0_en,
  input  [6:0]  W0_addr,
  input         W0_clk,
  input  [39:0] W0_data,
  input         W0_en
);
  wire [6:0] mem_0_0_iarp0;
  wire  mem_0_0_ickrp0;
  wire [39:0] mem_0_0_odoutp0;
  wire  mem_0_0_irenp0;
  wire [6:0] mem_0_0_iawp0;
  wire  mem_0_0_ickwp0;
  wire [39:0] mem_0_0_idinp0;
  wire  mem_0_0_iwenp0;
  wire  mem_0_0_ifuse;
  wire  mem_0_0_iclkbyp;
  wire  mem_0_0_imce;
  wire [1:0] mem_0_0_irmce;
  wire [3:0] mem_0_0_iwmce;
  wire [39:0] R0_data_0_0 = mem_0_0_odoutp0;
  wire [39:0] R0_data_0 = R0_data_0_0;
  ip224rfsbhpm1r1w128x40m1 mem_0_0 (
    .iarp0(mem_0_0_iarp0),
    .ickrp0(mem_0_0_ickrp0),
    .odoutp0(mem_0_0_odoutp0),
    .irenp0(mem_0_0_irenp0),
    .iawp0(mem_0_0_iawp0),
    .ickwp0(mem_0_0_ickwp0),
    .idinp0(mem_0_0_idinp0),
    .iwenp0(mem_0_0_iwenp0),
    .ifuse(mem_0_0_ifuse),
    .iclkbyp(mem_0_0_iclkbyp),
    .imce(mem_0_0_imce),
    .irmce(mem_0_0_irmce),
    .iwmce(mem_0_0_iwmce)
  );
  assign R0_data = mem_0_0_odoutp0;
  assign mem_0_0_iarp0 = R0_addr;
  assign mem_0_0_ickrp0 = R0_clk;
  assign mem_0_0_irenp0 = R0_en;
  assign mem_0_0_iawp0 = W0_addr;
  assign mem_0_0_ickwp0 = W0_clk;
  assign mem_0_0_idinp0 = W0_data;
  assign mem_0_0_iwenp0 = W0_en;
  assign mem_0_0_ifuse = 1'h0;
  assign mem_0_0_iclkbyp = 1'h0;
  assign mem_0_0_imce = 1'h0;
  assign mem_0_0_irmce = 2'h0;
  assign mem_0_0_iwmce = 4'h0;
endmodule
module data_ext(
  input  [10:0] R0_addr,
  input         R0_clk,
  output [7:0]  R0_data,
  input         R0_en,
  input  [10:0] W0_addr,
  input         W0_clk,
  input  [7:0]  W0_data,
  input         W0_en,
  input  [3:0]  W0_mask
);
  wire [10:0] mem_0_0_iarp0;
  wire  mem_0_0_ickrp0;
  wire [7:0] mem_0_0_odoutp0;
  wire  mem_0_0_irenp0;
  wire [10:0] mem_0_0_iawp0;
  wire  mem_0_0_ickwp0;
  wire [7:0] mem_0_0_idinp0;
  wire  mem_0_0_iwenp0;
  wire [7:0] mem_0_0_ibwep0;
  wire  mem_0_0_ifuse;
  wire  mem_0_0_iclkbyp;
  wire  mem_0_0_imce;
  wire [1:0] mem_0_0_irmce;
  wire [3:0] mem_0_0_iwmce;
  wire [7:0] R0_data_0_0 = mem_0_0_odoutp0;
  wire [7:0] R0_data_0 = R0_data_0_0;
  wire  _GEN_0 = W0_mask[0];
  wire  _GEN_1 = W0_mask[0];
  wire  _GEN_2 = W0_mask[1];
  wire [1:0] _GEN_3 = {W0_mask[0],W0_mask[0]};
  wire  _GEN_4 = W0_mask[1];
  wire [2:0] _GEN_5 = {W0_mask[1],W0_mask[0],W0_mask[0]};
  wire  _GEN_6 = W0_mask[2];
  wire [3:0] _GEN_7 = {W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0]};
  wire  _GEN_8 = W0_mask[2];
  wire [4:0] _GEN_9 = {W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0]};
  wire  _GEN_10 = W0_mask[3];
  wire [5:0] _GEN_11 = {W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0]};
  wire  _GEN_12 = W0_mask[3];
  wire [6:0] _GEN_13 = {W0_mask[3],W0_mask[2],W0_mask[2],W0_mask[1],W0_mask[1],W0_mask[0],W0_mask[0]};
  ip224rfsbhpm1r1w2048x8be8m4 mem_0_0 (
    .iarp0(mem_0_0_iarp0),
    .ickrp0(mem_0_0_ickrp0),
    .odoutp0(mem_0_0_odoutp0),
    .irenp0(mem_0_0_irenp0),
    .iawp0(mem_0_0_iawp0),
    .ickwp0(mem_0_0_ickwp0),
    .idinp0(mem_0_0_idinp0),
    .iwenp0(mem_0_0_iwenp0),
    .ibwep0(mem_0_0_ibwep0),
    .ifuse(mem_0_0_ifuse),
    .iclkbyp(mem_0_0_iclkbyp),
    .imce(mem_0_0_imce),
    .irmce(mem_0_0_irmce),
    .iwmce(mem_0_0_iwmce)
  );
  assign R0_data = mem_0_0_odoutp0;
  assign mem_0_0_iarp0 = R0_addr;
  assign mem_0_0_ickrp0 = R0_clk;
  assign mem_0_0_irenp0 = R0_en;
  assign mem_0_0_iawp0 = W0_addr;
  assign mem_0_0_ickwp0 = W0_clk;
  assign mem_0_0_idinp0 = W0_data;
  assign mem_0_0_iwenp0 = W0_en;
  assign mem_0_0_ibwep0 = {W0_mask[3],_GEN_13};
  assign mem_0_0_ifuse = 1'h0;
  assign mem_0_0_iclkbyp = 1'h0;
  assign mem_0_0_imce = 1'h0;
  assign mem_0_0_irmce = 2'h0;
  assign mem_0_0_iwmce = 4'h0;
endmodule
module meta_0_0_ext(
  input  [3:0]  R0_addr,
  input         R0_clk,
  output [49:0] R0_data,
  input         R0_en,
  input  [3:0]  W0_addr,
  input         W0_clk,
  input  [49:0] W0_data,
  input         W0_en
);
  wire [3:0] mem_0_0_iarp0;
  wire  mem_0_0_ickrp0;
  wire [63:0] mem_0_0_odoutp0;
  wire  mem_0_0_irenp0;
  wire [3:0] mem_0_0_iawp0;
  wire  mem_0_0_ickwp0;
  wire [63:0] mem_0_0_idinp0;
  wire  mem_0_0_iwenp0;
  wire  mem_0_0_ifuse;
  wire  mem_0_0_iclkbyp;
  wire  mem_0_0_imce;
  wire [1:0] mem_0_0_irmce;
  wire [3:0] mem_0_0_iwmce;
  wire [49:0] R0_data_0_0 = mem_0_0_odoutp0[49:0];
  wire [49:0] R0_data_0 = R0_data_0_0;
  ip224rfsbhpm1r1w16x64m2 mem_0_0 (
    .iarp0(mem_0_0_iarp0),
    .ickrp0(mem_0_0_ickrp0),
    .odoutp0(mem_0_0_odoutp0),
    .irenp0(mem_0_0_irenp0),
    .iawp0(mem_0_0_iawp0),
    .ickwp0(mem_0_0_ickwp0),
    .idinp0(mem_0_0_idinp0),
    .iwenp0(mem_0_0_iwenp0),
    .ifuse(mem_0_0_ifuse),
    .iclkbyp(mem_0_0_iclkbyp),
    .imce(mem_0_0_imce),
    .irmce(mem_0_0_irmce),
    .iwmce(mem_0_0_iwmce)
  );
  assign R0_data = mem_0_0_odoutp0[49:0];
  assign mem_0_0_iarp0 = R0_addr;
  assign mem_0_0_ickrp0 = R0_clk;
  assign mem_0_0_irenp0 = R0_en;
  assign mem_0_0_iawp0 = W0_addr;
  assign mem_0_0_ickwp0 = W0_clk;
  assign mem_0_0_idinp0 = {{14'd0}, W0_data};
  assign mem_0_0_iwenp0 = W0_en;
  assign mem_0_0_ifuse = 1'h0;
  assign mem_0_0_iclkbyp = 1'h0;
  assign mem_0_0_imce = 1'h0;
  assign mem_0_0_irmce = 2'h0;
  assign mem_0_0_iwmce = 4'h0;
endmodule
module ghist_0_ext(
  input  [3:0]  R0_addr,
  input         R0_clk,
  output [23:0] R0_data,
  input         R0_en,
  input  [3:0]  W0_addr,
  input         W0_clk,
  input  [23:0] W0_data,
  input         W0_en
);
  wire [3:0] mem_0_0_iarp0;
  wire  mem_0_0_ickrp0;
  wire [7:0] mem_0_0_odoutp0;
  wire  mem_0_0_irenp0;
  wire [3:0] mem_0_0_iawp0;
  wire  mem_0_0_ickwp0;
  wire [7:0] mem_0_0_idinp0;
  wire  mem_0_0_iwenp0;
  wire  mem_0_0_ifuse;
  wire  mem_0_0_iclkbyp;
  wire  mem_0_0_imce;
  wire [1:0] mem_0_0_irmce;
  wire [3:0] mem_0_0_iwmce;
  wire [3:0] mem_0_1_iarp0;
  wire  mem_0_1_ickrp0;
  wire [7:0] mem_0_1_odoutp0;
  wire  mem_0_1_irenp0;
  wire [3:0] mem_0_1_iawp0;
  wire  mem_0_1_ickwp0;
  wire [7:0] mem_0_1_idinp0;
  wire  mem_0_1_iwenp0;
  wire  mem_0_1_ifuse;
  wire  mem_0_1_iclkbyp;
  wire  mem_0_1_imce;
  wire [1:0] mem_0_1_irmce;
  wire [3:0] mem_0_1_iwmce;
  wire [3:0] mem_0_2_iarp0;
  wire  mem_0_2_ickrp0;
  wire [7:0] mem_0_2_odoutp0;
  wire  mem_0_2_irenp0;
  wire [3:0] mem_0_2_iawp0;
  wire  mem_0_2_ickwp0;
  wire [7:0] mem_0_2_idinp0;
  wire  mem_0_2_iwenp0;
  wire  mem_0_2_ifuse;
  wire  mem_0_2_iclkbyp;
  wire  mem_0_2_imce;
  wire [1:0] mem_0_2_irmce;
  wire [3:0] mem_0_2_iwmce;
  wire [7:0] R0_data_0_0 = mem_0_0_odoutp0;
  wire [7:0] R0_data_0_1 = mem_0_1_odoutp0;
  wire [7:0] R0_data_0_2 = mem_0_2_odoutp0;
  wire [15:0] _GEN_0 = {R0_data_0_1,R0_data_0_0};
  wire [23:0] R0_data_0 = {R0_data_0_2,R0_data_0_1,R0_data_0_0};
  wire [15:0] _GEN_1 = {R0_data_0_1,R0_data_0_0};
  ip224rfsbhpm1r1w16x8m1 mem_0_0 (
    .iarp0(mem_0_0_iarp0),
    .ickrp0(mem_0_0_ickrp0),
    .odoutp0(mem_0_0_odoutp0),
    .irenp0(mem_0_0_irenp0),
    .iawp0(mem_0_0_iawp0),
    .ickwp0(mem_0_0_ickwp0),
    .idinp0(mem_0_0_idinp0),
    .iwenp0(mem_0_0_iwenp0),
    .ifuse(mem_0_0_ifuse),
    .iclkbyp(mem_0_0_iclkbyp),
    .imce(mem_0_0_imce),
    .irmce(mem_0_0_irmce),
    .iwmce(mem_0_0_iwmce)
  );
  ip224rfsbhpm1r1w16x8m1 mem_0_1 (
    .iarp0(mem_0_1_iarp0),
    .ickrp0(mem_0_1_ickrp0),
    .odoutp0(mem_0_1_odoutp0),
    .irenp0(mem_0_1_irenp0),
    .iawp0(mem_0_1_iawp0),
    .ickwp0(mem_0_1_ickwp0),
    .idinp0(mem_0_1_idinp0),
    .iwenp0(mem_0_1_iwenp0),
    .ifuse(mem_0_1_ifuse),
    .iclkbyp(mem_0_1_iclkbyp),
    .imce(mem_0_1_imce),
    .irmce(mem_0_1_irmce),
    .iwmce(mem_0_1_iwmce)
  );
  ip224rfsbhpm1r1w16x8m1 mem_0_2 (
    .iarp0(mem_0_2_iarp0),
    .ickrp0(mem_0_2_ickrp0),
    .odoutp0(mem_0_2_odoutp0),
    .irenp0(mem_0_2_irenp0),
    .iawp0(mem_0_2_iawp0),
    .ickwp0(mem_0_2_ickwp0),
    .idinp0(mem_0_2_idinp0),
    .iwenp0(mem_0_2_iwenp0),
    .ifuse(mem_0_2_ifuse),
    .iclkbyp(mem_0_2_iclkbyp),
    .imce(mem_0_2_imce),
    .irmce(mem_0_2_irmce),
    .iwmce(mem_0_2_iwmce)
  );
  assign R0_data = {R0_data_0_2,_GEN_0};
  assign mem_0_0_iarp0 = R0_addr;
  assign mem_0_0_ickrp0 = R0_clk;
  assign mem_0_0_irenp0 = R0_en;
  assign mem_0_0_iawp0 = W0_addr;
  assign mem_0_0_ickwp0 = W0_clk;
  assign mem_0_0_idinp0 = W0_data[7:0];
  assign mem_0_0_iwenp0 = W0_en;
  assign mem_0_0_ifuse = 1'h0;
  assign mem_0_0_iclkbyp = 1'h0;
  assign mem_0_0_imce = 1'h0;
  assign mem_0_0_irmce = 2'h0;
  assign mem_0_0_iwmce = 4'h0;
  assign mem_0_1_iarp0 = R0_addr;
  assign mem_0_1_ickrp0 = R0_clk;
  assign mem_0_1_irenp0 = R0_en;
  assign mem_0_1_iawp0 = W0_addr;
  assign mem_0_1_ickwp0 = W0_clk;
  assign mem_0_1_idinp0 = W0_data[15:8];
  assign mem_0_1_iwenp0 = W0_en;
  assign mem_0_1_ifuse = 1'h0;
  assign mem_0_1_iclkbyp = 1'h0;
  assign mem_0_1_imce = 1'h0;
  assign mem_0_1_irmce = 2'h0;
  assign mem_0_1_iwmce = 4'h0;
  assign mem_0_2_iarp0 = R0_addr;
  assign mem_0_2_ickrp0 = R0_clk;
  assign mem_0_2_irenp0 = R0_en;
  assign mem_0_2_iawp0 = W0_addr;
  assign mem_0_2_ickwp0 = W0_clk;
  assign mem_0_2_idinp0 = W0_data[23:16];
  assign mem_0_2_iwenp0 = W0_en;
  assign mem_0_2_ifuse = 1'h0;
  assign mem_0_2_iclkbyp = 1'h0;
  assign mem_0_2_imce = 1'h0;
  assign mem_0_2_irmce = 2'h0;
  assign mem_0_2_iwmce = 4'h0;
endmodule
module rob_debug_inst_mem_0_ext(
  input  [4:0]  R0_addr,
  input         R0_clk,
  output [31:0] R0_data,
  input         R0_en,
  input  [4:0]  W0_addr,
  input         W0_clk,
  input  [31:0] W0_data,
  input         W0_en
);
  wire [4:0] mem_0_0_iarp0;
  wire  mem_0_0_ickrp0;
  wire [31:0] mem_0_0_odoutp0;
  wire  mem_0_0_irenp0;
  wire [4:0] mem_0_0_iawp0;
  wire  mem_0_0_ickwp0;
  wire [31:0] mem_0_0_idinp0;
  wire  mem_0_0_iwenp0;
  wire  mem_0_0_ifuse;
  wire  mem_0_0_iclkbyp;
  wire  mem_0_0_imce;
  wire [1:0] mem_0_0_irmce;
  wire [3:0] mem_0_0_iwmce;
  wire [31:0] R0_data_0_0 = mem_0_0_odoutp0;
  wire [31:0] R0_data_0 = R0_data_0_0;
  ip224rfsbhpm1r1w32x32m1 mem_0_0 (
    .iarp0(mem_0_0_iarp0),
    .ickrp0(mem_0_0_ickrp0),
    .odoutp0(mem_0_0_odoutp0),
    .irenp0(mem_0_0_irenp0),
    .iawp0(mem_0_0_iawp0),
    .ickwp0(mem_0_0_ickwp0),
    .idinp0(mem_0_0_idinp0),
    .iwenp0(mem_0_0_iwenp0),
    .ifuse(mem_0_0_ifuse),
    .iclkbyp(mem_0_0_iclkbyp),
    .imce(mem_0_0_imce),
    .irmce(mem_0_0_irmce),
    .iwmce(mem_0_0_iwmce)
  );
  assign R0_data = mem_0_0_odoutp0;
  assign mem_0_0_iarp0 = R0_addr;
  assign mem_0_0_ickrp0 = R0_clk;
  assign mem_0_0_irenp0 = R0_en;
  assign mem_0_0_iawp0 = W0_addr;
  assign mem_0_0_ickwp0 = W0_clk;
  assign mem_0_0_idinp0 = W0_data;
  assign mem_0_0_iwenp0 = W0_en;
  assign mem_0_0_ifuse = 1'h0;
  assign mem_0_0_iclkbyp = 1'h0;
  assign mem_0_0_imce = 1'h0;
  assign mem_0_0_irmce = 2'h0;
  assign mem_0_0_iwmce = 4'h0;
endmodule
