module signaltap (
		input  wire [63:0] acq_data_in,    //     tap.acq_data_in
		input  wire [31:0] acq_trigger_in, //        .acq_trigger_in
		input  wire        acq_clk         // acq_clk.clk
	);
endmodule

