module ring_terminator_n1 (
);

endmodule
